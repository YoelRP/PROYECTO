module counter(out, clk, reset);

  

endmodule // counter