////////////////////////////////////////////////////////////////////////////////
// Copyright (C) 1999-2008 Easics NV.
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//
// Purpose : synthesizable CRC function
//   * polynomial: x^16 + x^12 + x^5 + 1
//   * data width: 1024
//
// Info : tools@easics.be
//        http://www.easics.com
////////////////////////////////////////////////////////////////////////////////
module CRC16_D1024(
  nextCRC16_D1024,
  Data,
  crc
  );

  output reg  [15:0] nextCRC16_D1024;

    input wire [1023:0] Data;
    input wire [15:0] crc;
    reg [1023:0] d;
    reg [15:0] c;
    reg [15:0] newcrc;
  always @ (*) 
  begin
    d = Data;
    c = crc;

    newcrc[0] = d[1023] ^ d[1021] ^ d[1020] ^ d[1017] ^ d[1016] ^ d[1014] ^ d[1012] ^ d[1011] ^ d[1006] ^ d[1002] ^ d[999] ^ d[998] ^ d[997] ^ d[996] ^ d[995] ^ d[993] ^ d[992] ^ d[991] ^ d[990] ^ d[988] ^ d[986] ^ d[984] ^ d[983] ^ d[982] ^ d[981] ^ d[979] ^ d[976] ^ d[975] ^ d[974] ^ d[970] ^ d[968] ^ d[966] ^ d[964] ^ d[963] ^ d[962] ^ d[961] ^ d[960] ^ d[958] ^ d[957] ^ d[955] ^ d[953] ^ d[952] ^ d[951] ^ d[950] ^ d[949] ^ d[948] ^ d[946] ^ d[945] ^ d[942] ^ d[941] ^ d[938] ^ d[937] ^ d[936] ^ d[935] ^ d[933] ^ d[931] ^ d[930] ^ d[928] ^ d[926] ^ d[925] ^ d[924] ^ d[922] ^ d[921] ^ d[919] ^ d[918] ^ d[915] ^ d[914] ^ d[910] ^ d[909] ^ d[908] ^ d[907] ^ d[904] ^ d[903] ^ d[902] ^ d[898] ^ d[896] ^ d[895] ^ d[894] ^ d[891] ^ d[889] ^ d[888] ^ d[887] ^ d[886] ^ d[882] ^ d[881] ^ d[880] ^ d[878] ^ d[875] ^ d[874] ^ d[872] ^ d[871] ^ d[870] ^ d[868] ^ d[867] ^ d[866] ^ d[864] ^ d[862] ^ d[861] ^ d[860] ^ d[859] ^ d[857] ^ d[856] ^ d[855] ^ d[854] ^ d[852] ^ d[850] ^ d[846] ^ d[845] ^ d[842] ^ d[840] ^ d[839] ^ d[837] ^ d[836] ^ d[835] ^ d[834] ^ d[833] ^ d[832] ^ d[831] ^ d[830] ^ d[822] ^ d[816] ^ d[815] ^ d[814] ^ d[811] ^ d[809] ^ d[803] ^ d[802] ^ d[800] ^ d[793] ^ d[791] ^ d[790] ^ d[787] ^ d[785] ^ d[784] ^ d[782] ^ d[781] ^ d[780] ^ d[778] ^ d[776] ^ d[775] ^ d[774] ^ d[772] ^ d[769] ^ d[767] ^ d[765] ^ d[764] ^ d[763] ^ d[762] ^ d[760] ^ d[756] ^ d[752] ^ d[751] ^ d[750] ^ d[749] ^ d[745] ^ d[744] ^ d[740] ^ d[738] ^ d[737] ^ d[736] ^ d[734] ^ d[733] ^ d[731] ^ d[728] ^ d[725] ^ d[723] ^ d[719] ^ d[717] ^ d[716] ^ d[715] ^ d[714] ^ d[713] ^ d[710] ^ d[708] ^ d[704] ^ d[703] ^ d[702] ^ d[700] ^ d[698] ^ d[696] ^ d[695] ^ d[694] ^ d[693] ^ d[689] ^ d[688] ^ d[687] ^ d[684] ^ d[682] ^ d[681] ^ d[680] ^ d[678] ^ d[677] ^ d[672] ^ d[671] ^ d[670] ^ d[669] ^ d[667] ^ d[666] ^ d[665] ^ d[659] ^ d[658] ^ d[657] ^ d[656] ^ d[654] ^ d[653] ^ d[652] ^ d[650] ^ d[648] ^ d[646] ^ d[644] ^ d[641] ^ d[639] ^ d[637] ^ d[636] ^ d[634] ^ d[632] ^ d[631] ^ d[630] ^ d[628] ^ d[626] ^ d[625] ^ d[624] ^ d[622] ^ d[620] ^ d[617] ^ d[613] ^ d[612] ^ d[609] ^ d[608] ^ d[607] ^ d[606] ^ d[605] ^ d[603] ^ d[602] ^ d[601] ^ d[598] ^ d[597] ^ d[596] ^ d[595] ^ d[594] ^ d[593] ^ d[591] ^ d[590] ^ d[589] ^ d[588] ^ d[587] ^ d[586] ^ d[585] ^ d[582] ^ d[581] ^ d[577] ^ d[571] ^ d[561] ^ d[559] ^ d[556] ^ d[555] ^ d[554] ^ d[551] ^ d[550] ^ d[547] ^ d[546] ^ d[544] ^ d[541] ^ d[540] ^ d[539] ^ d[536] ^ d[535] ^ d[534] ^ d[532] ^ d[525] ^ d[522] ^ d[520] ^ d[519] ^ d[518] ^ d[517] ^ d[516] ^ d[515] ^ d[514] ^ d[512] ^ d[511] ^ d[508] ^ d[506] ^ d[505] ^ d[503] ^ d[500] ^ d[494] ^ d[493] ^ d[492] ^ d[491] ^ d[490] ^ d[486] ^ d[485] ^ d[484] ^ d[482] ^ d[476] ^ d[475] ^ d[473] ^ d[472] ^ d[471] ^ d[470] ^ d[469] ^ d[467] ^ d[465] ^ d[463] ^ d[462] ^ d[461] ^ d[460] ^ d[457] ^ d[455] ^ d[454] ^ d[452] ^ d[449] ^ d[448] ^ d[446] ^ d[442] ^ d[440] ^ d[439] ^ d[438] ^ d[435] ^ d[432] ^ d[430] ^ d[428] ^ d[425] ^ d[424] ^ d[423] ^ d[422] ^ d[417] ^ d[414] ^ d[413] ^ d[412] ^ d[411] ^ d[410] ^ d[402] ^ d[400] ^ d[399] ^ d[396] ^ d[391] ^ d[390] ^ d[388] ^ d[387] ^ d[385] ^ d[382] ^ d[379] ^ d[378] ^ d[377] ^ d[376] ^ d[370] ^ d[369] ^ d[367] ^ d[363] ^ d[361] ^ d[360] ^ d[357] ^ d[356] ^ d[354] ^ d[353] ^ d[352] ^ d[351] ^ d[346] ^ d[342] ^ d[341] ^ d[339] ^ d[338] ^ d[335] ^ d[333] ^ d[330] ^ d[329] ^ d[328] ^ d[327] ^ d[324] ^ d[323] ^ d[321] ^ d[315] ^ d[314] ^ d[313] ^ d[310] ^ d[307] ^ d[303] ^ d[301] ^ d[299] ^ d[298] ^ d[297] ^ d[296] ^ d[295] ^ d[293] ^ d[292] ^ d[291] ^ d[290] ^ d[289] ^ d[288] ^ d[287] ^ d[285] ^ d[283] ^ d[280] ^ d[275] ^ d[274] ^ d[272] ^ d[270] ^ d[268] ^ d[265] ^ d[264] ^ d[262] ^ d[257] ^ d[254] ^ d[253] ^ d[252] ^ d[250] ^ d[247] ^ d[246] ^ d[241] ^ d[240] ^ d[237] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[222] ^ d[219] ^ d[214] ^ d[212] ^ d[207] ^ d[206] ^ d[203] ^ d[201] ^ d[200] ^ d[194] ^ d[190] ^ d[188] ^ d[187] ^ d[184] ^ d[183] ^ d[179] ^ d[178] ^ d[176] ^ d[175] ^ d[173] ^ d[171] ^ d[170] ^ d[165] ^ d[164] ^ d[162] ^ d[161] ^ d[159] ^ d[158] ^ d[156] ^ d[155] ^ d[152] ^ d[151] ^ d[148] ^ d[146] ^ d[145] ^ d[144] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[132] ^ d[127] ^ d[123] ^ d[121] ^ d[118] ^ d[115] ^ d[113] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[104] ^ d[98] ^ d[96] ^ d[95] ^ d[88] ^ d[86] ^ d[84] ^ d[82] ^ d[81] ^ d[80] ^ d[77] ^ d[75] ^ d[74] ^ d[72] ^ d[70] ^ d[67] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[58] ^ d[56] ^ d[55] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[42] ^ d[35] ^ d[33] ^ d[32] ^ d[28] ^ d[27] ^ d[26] ^ d[22] ^ d[20] ^ d[19] ^ d[12] ^ d[11] ^ d[8] ^ d[4] ^ d[0] ^ c[3] ^ c[4] ^ c[6] ^ c[8] ^ c[9] ^ c[12] ^ c[13] ^ c[15];
    newcrc[1] = d[1022] ^ d[1021] ^ d[1018] ^ d[1017] ^ d[1015] ^ d[1013] ^ d[1012] ^ d[1007] ^ d[1003] ^ d[1000] ^ d[999] ^ d[998] ^ d[997] ^ d[996] ^ d[994] ^ d[993] ^ d[992] ^ d[991] ^ d[989] ^ d[987] ^ d[985] ^ d[984] ^ d[983] ^ d[982] ^ d[980] ^ d[977] ^ d[976] ^ d[975] ^ d[971] ^ d[969] ^ d[967] ^ d[965] ^ d[964] ^ d[963] ^ d[962] ^ d[961] ^ d[959] ^ d[958] ^ d[956] ^ d[954] ^ d[953] ^ d[952] ^ d[951] ^ d[950] ^ d[949] ^ d[947] ^ d[946] ^ d[943] ^ d[942] ^ d[939] ^ d[938] ^ d[937] ^ d[936] ^ d[934] ^ d[932] ^ d[931] ^ d[929] ^ d[927] ^ d[926] ^ d[925] ^ d[923] ^ d[922] ^ d[920] ^ d[919] ^ d[916] ^ d[915] ^ d[911] ^ d[910] ^ d[909] ^ d[908] ^ d[905] ^ d[904] ^ d[903] ^ d[899] ^ d[897] ^ d[896] ^ d[895] ^ d[892] ^ d[890] ^ d[889] ^ d[888] ^ d[887] ^ d[883] ^ d[882] ^ d[881] ^ d[879] ^ d[876] ^ d[875] ^ d[873] ^ d[872] ^ d[871] ^ d[869] ^ d[868] ^ d[867] ^ d[865] ^ d[863] ^ d[862] ^ d[861] ^ d[860] ^ d[858] ^ d[857] ^ d[856] ^ d[855] ^ d[853] ^ d[851] ^ d[847] ^ d[846] ^ d[843] ^ d[841] ^ d[840] ^ d[838] ^ d[837] ^ d[836] ^ d[835] ^ d[834] ^ d[833] ^ d[832] ^ d[831] ^ d[823] ^ d[817] ^ d[816] ^ d[815] ^ d[812] ^ d[810] ^ d[804] ^ d[803] ^ d[801] ^ d[794] ^ d[792] ^ d[791] ^ d[788] ^ d[786] ^ d[785] ^ d[783] ^ d[782] ^ d[781] ^ d[779] ^ d[777] ^ d[776] ^ d[775] ^ d[773] ^ d[770] ^ d[768] ^ d[766] ^ d[765] ^ d[764] ^ d[763] ^ d[761] ^ d[757] ^ d[753] ^ d[752] ^ d[751] ^ d[750] ^ d[746] ^ d[745] ^ d[741] ^ d[739] ^ d[738] ^ d[737] ^ d[735] ^ d[734] ^ d[732] ^ d[729] ^ d[726] ^ d[724] ^ d[720] ^ d[718] ^ d[717] ^ d[716] ^ d[715] ^ d[714] ^ d[711] ^ d[709] ^ d[705] ^ d[704] ^ d[703] ^ d[701] ^ d[699] ^ d[697] ^ d[696] ^ d[695] ^ d[694] ^ d[690] ^ d[689] ^ d[688] ^ d[685] ^ d[683] ^ d[682] ^ d[681] ^ d[679] ^ d[678] ^ d[673] ^ d[672] ^ d[671] ^ d[670] ^ d[668] ^ d[667] ^ d[666] ^ d[660] ^ d[659] ^ d[658] ^ d[657] ^ d[655] ^ d[654] ^ d[653] ^ d[651] ^ d[649] ^ d[647] ^ d[645] ^ d[642] ^ d[640] ^ d[638] ^ d[637] ^ d[635] ^ d[633] ^ d[632] ^ d[631] ^ d[629] ^ d[627] ^ d[626] ^ d[625] ^ d[623] ^ d[621] ^ d[618] ^ d[614] ^ d[613] ^ d[610] ^ d[609] ^ d[608] ^ d[607] ^ d[606] ^ d[604] ^ d[603] ^ d[602] ^ d[599] ^ d[598] ^ d[597] ^ d[596] ^ d[595] ^ d[594] ^ d[592] ^ d[591] ^ d[590] ^ d[589] ^ d[588] ^ d[587] ^ d[586] ^ d[583] ^ d[582] ^ d[578] ^ d[572] ^ d[562] ^ d[560] ^ d[557] ^ d[556] ^ d[555] ^ d[552] ^ d[551] ^ d[548] ^ d[547] ^ d[545] ^ d[542] ^ d[541] ^ d[540] ^ d[537] ^ d[536] ^ d[535] ^ d[533] ^ d[526] ^ d[523] ^ d[521] ^ d[520] ^ d[519] ^ d[518] ^ d[517] ^ d[516] ^ d[515] ^ d[513] ^ d[512] ^ d[509] ^ d[507] ^ d[506] ^ d[504] ^ d[501] ^ d[495] ^ d[494] ^ d[493] ^ d[492] ^ d[491] ^ d[487] ^ d[486] ^ d[485] ^ d[483] ^ d[477] ^ d[476] ^ d[474] ^ d[473] ^ d[472] ^ d[471] ^ d[470] ^ d[468] ^ d[466] ^ d[464] ^ d[463] ^ d[462] ^ d[461] ^ d[458] ^ d[456] ^ d[455] ^ d[453] ^ d[450] ^ d[449] ^ d[447] ^ d[443] ^ d[441] ^ d[440] ^ d[439] ^ d[436] ^ d[433] ^ d[431] ^ d[429] ^ d[426] ^ d[425] ^ d[424] ^ d[423] ^ d[418] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[411] ^ d[403] ^ d[401] ^ d[400] ^ d[397] ^ d[392] ^ d[391] ^ d[389] ^ d[388] ^ d[386] ^ d[383] ^ d[380] ^ d[379] ^ d[378] ^ d[377] ^ d[371] ^ d[370] ^ d[368] ^ d[364] ^ d[362] ^ d[361] ^ d[358] ^ d[357] ^ d[355] ^ d[354] ^ d[353] ^ d[352] ^ d[347] ^ d[343] ^ d[342] ^ d[340] ^ d[339] ^ d[336] ^ d[334] ^ d[331] ^ d[330] ^ d[329] ^ d[328] ^ d[325] ^ d[324] ^ d[322] ^ d[316] ^ d[315] ^ d[314] ^ d[311] ^ d[308] ^ d[304] ^ d[302] ^ d[300] ^ d[299] ^ d[298] ^ d[297] ^ d[296] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[290] ^ d[289] ^ d[288] ^ d[286] ^ d[284] ^ d[281] ^ d[276] ^ d[275] ^ d[273] ^ d[271] ^ d[269] ^ d[266] ^ d[265] ^ d[263] ^ d[258] ^ d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[248] ^ d[247] ^ d[242] ^ d[241] ^ d[238] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[224] ^ d[223] ^ d[220] ^ d[215] ^ d[213] ^ d[208] ^ d[207] ^ d[204] ^ d[202] ^ d[201] ^ d[195] ^ d[191] ^ d[189] ^ d[188] ^ d[185] ^ d[184] ^ d[180] ^ d[179] ^ d[177] ^ d[176] ^ d[174] ^ d[172] ^ d[171] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[160] ^ d[159] ^ d[157] ^ d[156] ^ d[153] ^ d[152] ^ d[149] ^ d[147] ^ d[146] ^ d[145] ^ d[144] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[133] ^ d[128] ^ d[124] ^ d[122] ^ d[119] ^ d[116] ^ d[114] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[99] ^ d[97] ^ d[96] ^ d[89] ^ d[87] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[78] ^ d[76] ^ d[75] ^ d[73] ^ d[71] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[64] ^ d[59] ^ d[57] ^ d[56] ^ d[53] ^ d[52] ^ d[50] ^ d[49] ^ d[43] ^ d[36] ^ d[34] ^ d[33] ^ d[29] ^ d[28] ^ d[27] ^ d[23] ^ d[21] ^ d[20] ^ d[13] ^ d[12] ^ d[9] ^ d[5] ^ d[1] ^ c[4] ^ c[5] ^ c[7] ^ c[9] ^ c[10] ^ c[13] ^ c[14];
    newcrc[2] = d[1023] ^ d[1022] ^ d[1019] ^ d[1018] ^ d[1016] ^ d[1014] ^ d[1013] ^ d[1008] ^ d[1004] ^ d[1001] ^ d[1000] ^ d[999] ^ d[998] ^ d[997] ^ d[995] ^ d[994] ^ d[993] ^ d[992] ^ d[990] ^ d[988] ^ d[986] ^ d[985] ^ d[984] ^ d[983] ^ d[981] ^ d[978] ^ d[977] ^ d[976] ^ d[972] ^ d[970] ^ d[968] ^ d[966] ^ d[965] ^ d[964] ^ d[963] ^ d[962] ^ d[960] ^ d[959] ^ d[957] ^ d[955] ^ d[954] ^ d[953] ^ d[952] ^ d[951] ^ d[950] ^ d[948] ^ d[947] ^ d[944] ^ d[943] ^ d[940] ^ d[939] ^ d[938] ^ d[937] ^ d[935] ^ d[933] ^ d[932] ^ d[930] ^ d[928] ^ d[927] ^ d[926] ^ d[924] ^ d[923] ^ d[921] ^ d[920] ^ d[917] ^ d[916] ^ d[912] ^ d[911] ^ d[910] ^ d[909] ^ d[906] ^ d[905] ^ d[904] ^ d[900] ^ d[898] ^ d[897] ^ d[896] ^ d[893] ^ d[891] ^ d[890] ^ d[889] ^ d[888] ^ d[884] ^ d[883] ^ d[882] ^ d[880] ^ d[877] ^ d[876] ^ d[874] ^ d[873] ^ d[872] ^ d[870] ^ d[869] ^ d[868] ^ d[866] ^ d[864] ^ d[863] ^ d[862] ^ d[861] ^ d[859] ^ d[858] ^ d[857] ^ d[856] ^ d[854] ^ d[852] ^ d[848] ^ d[847] ^ d[844] ^ d[842] ^ d[841] ^ d[839] ^ d[838] ^ d[837] ^ d[836] ^ d[835] ^ d[834] ^ d[833] ^ d[832] ^ d[824] ^ d[818] ^ d[817] ^ d[816] ^ d[813] ^ d[811] ^ d[805] ^ d[804] ^ d[802] ^ d[795] ^ d[793] ^ d[792] ^ d[789] ^ d[787] ^ d[786] ^ d[784] ^ d[783] ^ d[782] ^ d[780] ^ d[778] ^ d[777] ^ d[776] ^ d[774] ^ d[771] ^ d[769] ^ d[767] ^ d[766] ^ d[765] ^ d[764] ^ d[762] ^ d[758] ^ d[754] ^ d[753] ^ d[752] ^ d[751] ^ d[747] ^ d[746] ^ d[742] ^ d[740] ^ d[739] ^ d[738] ^ d[736] ^ d[735] ^ d[733] ^ d[730] ^ d[727] ^ d[725] ^ d[721] ^ d[719] ^ d[718] ^ d[717] ^ d[716] ^ d[715] ^ d[712] ^ d[710] ^ d[706] ^ d[705] ^ d[704] ^ d[702] ^ d[700] ^ d[698] ^ d[697] ^ d[696] ^ d[695] ^ d[691] ^ d[690] ^ d[689] ^ d[686] ^ d[684] ^ d[683] ^ d[682] ^ d[680] ^ d[679] ^ d[674] ^ d[673] ^ d[672] ^ d[671] ^ d[669] ^ d[668] ^ d[667] ^ d[661] ^ d[660] ^ d[659] ^ d[658] ^ d[656] ^ d[655] ^ d[654] ^ d[652] ^ d[650] ^ d[648] ^ d[646] ^ d[643] ^ d[641] ^ d[639] ^ d[638] ^ d[636] ^ d[634] ^ d[633] ^ d[632] ^ d[630] ^ d[628] ^ d[627] ^ d[626] ^ d[624] ^ d[622] ^ d[619] ^ d[615] ^ d[614] ^ d[611] ^ d[610] ^ d[609] ^ d[608] ^ d[607] ^ d[605] ^ d[604] ^ d[603] ^ d[600] ^ d[599] ^ d[598] ^ d[597] ^ d[596] ^ d[595] ^ d[593] ^ d[592] ^ d[591] ^ d[590] ^ d[589] ^ d[588] ^ d[587] ^ d[584] ^ d[583] ^ d[579] ^ d[573] ^ d[563] ^ d[561] ^ d[558] ^ d[557] ^ d[556] ^ d[553] ^ d[552] ^ d[549] ^ d[548] ^ d[546] ^ d[543] ^ d[542] ^ d[541] ^ d[538] ^ d[537] ^ d[536] ^ d[534] ^ d[527] ^ d[524] ^ d[522] ^ d[521] ^ d[520] ^ d[519] ^ d[518] ^ d[517] ^ d[516] ^ d[514] ^ d[513] ^ d[510] ^ d[508] ^ d[507] ^ d[505] ^ d[502] ^ d[496] ^ d[495] ^ d[494] ^ d[493] ^ d[492] ^ d[488] ^ d[487] ^ d[486] ^ d[484] ^ d[478] ^ d[477] ^ d[475] ^ d[474] ^ d[473] ^ d[472] ^ d[471] ^ d[469] ^ d[467] ^ d[465] ^ d[464] ^ d[463] ^ d[462] ^ d[459] ^ d[457] ^ d[456] ^ d[454] ^ d[451] ^ d[450] ^ d[448] ^ d[444] ^ d[442] ^ d[441] ^ d[440] ^ d[437] ^ d[434] ^ d[432] ^ d[430] ^ d[427] ^ d[426] ^ d[425] ^ d[424] ^ d[419] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[404] ^ d[402] ^ d[401] ^ d[398] ^ d[393] ^ d[392] ^ d[390] ^ d[389] ^ d[387] ^ d[384] ^ d[381] ^ d[380] ^ d[379] ^ d[378] ^ d[372] ^ d[371] ^ d[369] ^ d[365] ^ d[363] ^ d[362] ^ d[359] ^ d[358] ^ d[356] ^ d[355] ^ d[354] ^ d[353] ^ d[348] ^ d[344] ^ d[343] ^ d[341] ^ d[340] ^ d[337] ^ d[335] ^ d[332] ^ d[331] ^ d[330] ^ d[329] ^ d[326] ^ d[325] ^ d[323] ^ d[317] ^ d[316] ^ d[315] ^ d[312] ^ d[309] ^ d[305] ^ d[303] ^ d[301] ^ d[300] ^ d[299] ^ d[298] ^ d[297] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[290] ^ d[289] ^ d[287] ^ d[285] ^ d[282] ^ d[277] ^ d[276] ^ d[274] ^ d[272] ^ d[270] ^ d[267] ^ d[266] ^ d[264] ^ d[259] ^ d[256] ^ d[255] ^ d[254] ^ d[252] ^ d[249] ^ d[248] ^ d[243] ^ d[242] ^ d[239] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[225] ^ d[224] ^ d[221] ^ d[216] ^ d[214] ^ d[209] ^ d[208] ^ d[205] ^ d[203] ^ d[202] ^ d[196] ^ d[192] ^ d[190] ^ d[189] ^ d[186] ^ d[185] ^ d[181] ^ d[180] ^ d[178] ^ d[177] ^ d[175] ^ d[173] ^ d[172] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[161] ^ d[160] ^ d[158] ^ d[157] ^ d[154] ^ d[153] ^ d[150] ^ d[148] ^ d[147] ^ d[146] ^ d[145] ^ d[144] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[134] ^ d[129] ^ d[125] ^ d[123] ^ d[120] ^ d[117] ^ d[115] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[100] ^ d[98] ^ d[97] ^ d[90] ^ d[88] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[79] ^ d[77] ^ d[76] ^ d[74] ^ d[72] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[60] ^ d[58] ^ d[57] ^ d[54] ^ d[53] ^ d[51] ^ d[50] ^ d[44] ^ d[37] ^ d[35] ^ d[34] ^ d[30] ^ d[29] ^ d[28] ^ d[24] ^ d[22] ^ d[21] ^ d[14] ^ d[13] ^ d[10] ^ d[6] ^ d[2] ^ c[0] ^ c[5] ^ c[6] ^ c[8] ^ c[10] ^ c[11] ^ c[14] ^ c[15];
    newcrc[3] = d[1023] ^ d[1020] ^ d[1019] ^ d[1017] ^ d[1015] ^ d[1014] ^ d[1009] ^ d[1005] ^ d[1002] ^ d[1001] ^ d[1000] ^ d[999] ^ d[998] ^ d[996] ^ d[995] ^ d[994] ^ d[993] ^ d[991] ^ d[989] ^ d[987] ^ d[986] ^ d[985] ^ d[984] ^ d[982] ^ d[979] ^ d[978] ^ d[977] ^ d[973] ^ d[971] ^ d[969] ^ d[967] ^ d[966] ^ d[965] ^ d[964] ^ d[963] ^ d[961] ^ d[960] ^ d[958] ^ d[956] ^ d[955] ^ d[954] ^ d[953] ^ d[952] ^ d[951] ^ d[949] ^ d[948] ^ d[945] ^ d[944] ^ d[941] ^ d[940] ^ d[939] ^ d[938] ^ d[936] ^ d[934] ^ d[933] ^ d[931] ^ d[929] ^ d[928] ^ d[927] ^ d[925] ^ d[924] ^ d[922] ^ d[921] ^ d[918] ^ d[917] ^ d[913] ^ d[912] ^ d[911] ^ d[910] ^ d[907] ^ d[906] ^ d[905] ^ d[901] ^ d[899] ^ d[898] ^ d[897] ^ d[894] ^ d[892] ^ d[891] ^ d[890] ^ d[889] ^ d[885] ^ d[884] ^ d[883] ^ d[881] ^ d[878] ^ d[877] ^ d[875] ^ d[874] ^ d[873] ^ d[871] ^ d[870] ^ d[869] ^ d[867] ^ d[865] ^ d[864] ^ d[863] ^ d[862] ^ d[860] ^ d[859] ^ d[858] ^ d[857] ^ d[855] ^ d[853] ^ d[849] ^ d[848] ^ d[845] ^ d[843] ^ d[842] ^ d[840] ^ d[839] ^ d[838] ^ d[837] ^ d[836] ^ d[835] ^ d[834] ^ d[833] ^ d[825] ^ d[819] ^ d[818] ^ d[817] ^ d[814] ^ d[812] ^ d[806] ^ d[805] ^ d[803] ^ d[796] ^ d[794] ^ d[793] ^ d[790] ^ d[788] ^ d[787] ^ d[785] ^ d[784] ^ d[783] ^ d[781] ^ d[779] ^ d[778] ^ d[777] ^ d[775] ^ d[772] ^ d[770] ^ d[768] ^ d[767] ^ d[766] ^ d[765] ^ d[763] ^ d[759] ^ d[755] ^ d[754] ^ d[753] ^ d[752] ^ d[748] ^ d[747] ^ d[743] ^ d[741] ^ d[740] ^ d[739] ^ d[737] ^ d[736] ^ d[734] ^ d[731] ^ d[728] ^ d[726] ^ d[722] ^ d[720] ^ d[719] ^ d[718] ^ d[717] ^ d[716] ^ d[713] ^ d[711] ^ d[707] ^ d[706] ^ d[705] ^ d[703] ^ d[701] ^ d[699] ^ d[698] ^ d[697] ^ d[696] ^ d[692] ^ d[691] ^ d[690] ^ d[687] ^ d[685] ^ d[684] ^ d[683] ^ d[681] ^ d[680] ^ d[675] ^ d[674] ^ d[673] ^ d[672] ^ d[670] ^ d[669] ^ d[668] ^ d[662] ^ d[661] ^ d[660] ^ d[659] ^ d[657] ^ d[656] ^ d[655] ^ d[653] ^ d[651] ^ d[649] ^ d[647] ^ d[644] ^ d[642] ^ d[640] ^ d[639] ^ d[637] ^ d[635] ^ d[634] ^ d[633] ^ d[631] ^ d[629] ^ d[628] ^ d[627] ^ d[625] ^ d[623] ^ d[620] ^ d[616] ^ d[615] ^ d[612] ^ d[611] ^ d[610] ^ d[609] ^ d[608] ^ d[606] ^ d[605] ^ d[604] ^ d[601] ^ d[600] ^ d[599] ^ d[598] ^ d[597] ^ d[596] ^ d[594] ^ d[593] ^ d[592] ^ d[591] ^ d[590] ^ d[589] ^ d[588] ^ d[585] ^ d[584] ^ d[580] ^ d[574] ^ d[564] ^ d[562] ^ d[559] ^ d[558] ^ d[557] ^ d[554] ^ d[553] ^ d[550] ^ d[549] ^ d[547] ^ d[544] ^ d[543] ^ d[542] ^ d[539] ^ d[538] ^ d[537] ^ d[535] ^ d[528] ^ d[525] ^ d[523] ^ d[522] ^ d[521] ^ d[520] ^ d[519] ^ d[518] ^ d[517] ^ d[515] ^ d[514] ^ d[511] ^ d[509] ^ d[508] ^ d[506] ^ d[503] ^ d[497] ^ d[496] ^ d[495] ^ d[494] ^ d[493] ^ d[489] ^ d[488] ^ d[487] ^ d[485] ^ d[479] ^ d[478] ^ d[476] ^ d[475] ^ d[474] ^ d[473] ^ d[472] ^ d[470] ^ d[468] ^ d[466] ^ d[465] ^ d[464] ^ d[463] ^ d[460] ^ d[458] ^ d[457] ^ d[455] ^ d[452] ^ d[451] ^ d[449] ^ d[445] ^ d[443] ^ d[442] ^ d[441] ^ d[438] ^ d[435] ^ d[433] ^ d[431] ^ d[428] ^ d[427] ^ d[426] ^ d[425] ^ d[420] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[405] ^ d[403] ^ d[402] ^ d[399] ^ d[394] ^ d[393] ^ d[391] ^ d[390] ^ d[388] ^ d[385] ^ d[382] ^ d[381] ^ d[380] ^ d[379] ^ d[373] ^ d[372] ^ d[370] ^ d[366] ^ d[364] ^ d[363] ^ d[360] ^ d[359] ^ d[357] ^ d[356] ^ d[355] ^ d[354] ^ d[349] ^ d[345] ^ d[344] ^ d[342] ^ d[341] ^ d[338] ^ d[336] ^ d[333] ^ d[332] ^ d[331] ^ d[330] ^ d[327] ^ d[326] ^ d[324] ^ d[318] ^ d[317] ^ d[316] ^ d[313] ^ d[310] ^ d[306] ^ d[304] ^ d[302] ^ d[301] ^ d[300] ^ d[299] ^ d[298] ^ d[296] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[290] ^ d[288] ^ d[286] ^ d[283] ^ d[278] ^ d[277] ^ d[275] ^ d[273] ^ d[271] ^ d[268] ^ d[267] ^ d[265] ^ d[260] ^ d[257] ^ d[256] ^ d[255] ^ d[253] ^ d[250] ^ d[249] ^ d[244] ^ d[243] ^ d[240] ^ d[235] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[226] ^ d[225] ^ d[222] ^ d[217] ^ d[215] ^ d[210] ^ d[209] ^ d[206] ^ d[204] ^ d[203] ^ d[197] ^ d[193] ^ d[191] ^ d[190] ^ d[187] ^ d[186] ^ d[182] ^ d[181] ^ d[179] ^ d[178] ^ d[176] ^ d[174] ^ d[173] ^ d[168] ^ d[167] ^ d[165] ^ d[164] ^ d[162] ^ d[161] ^ d[159] ^ d[158] ^ d[155] ^ d[154] ^ d[151] ^ d[149] ^ d[148] ^ d[147] ^ d[146] ^ d[145] ^ d[144] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[135] ^ d[130] ^ d[126] ^ d[124] ^ d[121] ^ d[118] ^ d[116] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[107] ^ d[101] ^ d[99] ^ d[98] ^ d[91] ^ d[89] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[80] ^ d[78] ^ d[77] ^ d[75] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[61] ^ d[59] ^ d[58] ^ d[55] ^ d[54] ^ d[52] ^ d[51] ^ d[45] ^ d[38] ^ d[36] ^ d[35] ^ d[31] ^ d[30] ^ d[29] ^ d[25] ^ d[23] ^ d[22] ^ d[15] ^ d[14] ^ d[11] ^ d[7] ^ d[3] ^ c[1] ^ c[6] ^ c[7] ^ c[9] ^ c[11] ^ c[12] ^ c[15];
    newcrc[4] = d[1021] ^ d[1020] ^ d[1018] ^ d[1016] ^ d[1015] ^ d[1010] ^ d[1006] ^ d[1003] ^ d[1002] ^ d[1001] ^ d[1000] ^ d[999] ^ d[997] ^ d[996] ^ d[995] ^ d[994] ^ d[992] ^ d[990] ^ d[988] ^ d[987] ^ d[986] ^ d[985] ^ d[983] ^ d[980] ^ d[979] ^ d[978] ^ d[974] ^ d[972] ^ d[970] ^ d[968] ^ d[967] ^ d[966] ^ d[965] ^ d[964] ^ d[962] ^ d[961] ^ d[959] ^ d[957] ^ d[956] ^ d[955] ^ d[954] ^ d[953] ^ d[952] ^ d[950] ^ d[949] ^ d[946] ^ d[945] ^ d[942] ^ d[941] ^ d[940] ^ d[939] ^ d[937] ^ d[935] ^ d[934] ^ d[932] ^ d[930] ^ d[929] ^ d[928] ^ d[926] ^ d[925] ^ d[923] ^ d[922] ^ d[919] ^ d[918] ^ d[914] ^ d[913] ^ d[912] ^ d[911] ^ d[908] ^ d[907] ^ d[906] ^ d[902] ^ d[900] ^ d[899] ^ d[898] ^ d[895] ^ d[893] ^ d[892] ^ d[891] ^ d[890] ^ d[886] ^ d[885] ^ d[884] ^ d[882] ^ d[879] ^ d[878] ^ d[876] ^ d[875] ^ d[874] ^ d[872] ^ d[871] ^ d[870] ^ d[868] ^ d[866] ^ d[865] ^ d[864] ^ d[863] ^ d[861] ^ d[860] ^ d[859] ^ d[858] ^ d[856] ^ d[854] ^ d[850] ^ d[849] ^ d[846] ^ d[844] ^ d[843] ^ d[841] ^ d[840] ^ d[839] ^ d[838] ^ d[837] ^ d[836] ^ d[835] ^ d[834] ^ d[826] ^ d[820] ^ d[819] ^ d[818] ^ d[815] ^ d[813] ^ d[807] ^ d[806] ^ d[804] ^ d[797] ^ d[795] ^ d[794] ^ d[791] ^ d[789] ^ d[788] ^ d[786] ^ d[785] ^ d[784] ^ d[782] ^ d[780] ^ d[779] ^ d[778] ^ d[776] ^ d[773] ^ d[771] ^ d[769] ^ d[768] ^ d[767] ^ d[766] ^ d[764] ^ d[760] ^ d[756] ^ d[755] ^ d[754] ^ d[753] ^ d[749] ^ d[748] ^ d[744] ^ d[742] ^ d[741] ^ d[740] ^ d[738] ^ d[737] ^ d[735] ^ d[732] ^ d[729] ^ d[727] ^ d[723] ^ d[721] ^ d[720] ^ d[719] ^ d[718] ^ d[717] ^ d[714] ^ d[712] ^ d[708] ^ d[707] ^ d[706] ^ d[704] ^ d[702] ^ d[700] ^ d[699] ^ d[698] ^ d[697] ^ d[693] ^ d[692] ^ d[691] ^ d[688] ^ d[686] ^ d[685] ^ d[684] ^ d[682] ^ d[681] ^ d[676] ^ d[675] ^ d[674] ^ d[673] ^ d[671] ^ d[670] ^ d[669] ^ d[663] ^ d[662] ^ d[661] ^ d[660] ^ d[658] ^ d[657] ^ d[656] ^ d[654] ^ d[652] ^ d[650] ^ d[648] ^ d[645] ^ d[643] ^ d[641] ^ d[640] ^ d[638] ^ d[636] ^ d[635] ^ d[634] ^ d[632] ^ d[630] ^ d[629] ^ d[628] ^ d[626] ^ d[624] ^ d[621] ^ d[617] ^ d[616] ^ d[613] ^ d[612] ^ d[611] ^ d[610] ^ d[609] ^ d[607] ^ d[606] ^ d[605] ^ d[602] ^ d[601] ^ d[600] ^ d[599] ^ d[598] ^ d[597] ^ d[595] ^ d[594] ^ d[593] ^ d[592] ^ d[591] ^ d[590] ^ d[589] ^ d[586] ^ d[585] ^ d[581] ^ d[575] ^ d[565] ^ d[563] ^ d[560] ^ d[559] ^ d[558] ^ d[555] ^ d[554] ^ d[551] ^ d[550] ^ d[548] ^ d[545] ^ d[544] ^ d[543] ^ d[540] ^ d[539] ^ d[538] ^ d[536] ^ d[529] ^ d[526] ^ d[524] ^ d[523] ^ d[522] ^ d[521] ^ d[520] ^ d[519] ^ d[518] ^ d[516] ^ d[515] ^ d[512] ^ d[510] ^ d[509] ^ d[507] ^ d[504] ^ d[498] ^ d[497] ^ d[496] ^ d[495] ^ d[494] ^ d[490] ^ d[489] ^ d[488] ^ d[486] ^ d[480] ^ d[479] ^ d[477] ^ d[476] ^ d[475] ^ d[474] ^ d[473] ^ d[471] ^ d[469] ^ d[467] ^ d[466] ^ d[465] ^ d[464] ^ d[461] ^ d[459] ^ d[458] ^ d[456] ^ d[453] ^ d[452] ^ d[450] ^ d[446] ^ d[444] ^ d[443] ^ d[442] ^ d[439] ^ d[436] ^ d[434] ^ d[432] ^ d[429] ^ d[428] ^ d[427] ^ d[426] ^ d[421] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[406] ^ d[404] ^ d[403] ^ d[400] ^ d[395] ^ d[394] ^ d[392] ^ d[391] ^ d[389] ^ d[386] ^ d[383] ^ d[382] ^ d[381] ^ d[380] ^ d[374] ^ d[373] ^ d[371] ^ d[367] ^ d[365] ^ d[364] ^ d[361] ^ d[360] ^ d[358] ^ d[357] ^ d[356] ^ d[355] ^ d[350] ^ d[346] ^ d[345] ^ d[343] ^ d[342] ^ d[339] ^ d[337] ^ d[334] ^ d[333] ^ d[332] ^ d[331] ^ d[328] ^ d[327] ^ d[325] ^ d[319] ^ d[318] ^ d[317] ^ d[314] ^ d[311] ^ d[307] ^ d[305] ^ d[303] ^ d[302] ^ d[301] ^ d[300] ^ d[299] ^ d[297] ^ d[296] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[289] ^ d[287] ^ d[284] ^ d[279] ^ d[278] ^ d[276] ^ d[274] ^ d[272] ^ d[269] ^ d[268] ^ d[266] ^ d[261] ^ d[258] ^ d[257] ^ d[256] ^ d[254] ^ d[251] ^ d[250] ^ d[245] ^ d[244] ^ d[241] ^ d[236] ^ d[235] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[227] ^ d[226] ^ d[223] ^ d[218] ^ d[216] ^ d[211] ^ d[210] ^ d[207] ^ d[205] ^ d[204] ^ d[198] ^ d[194] ^ d[192] ^ d[191] ^ d[188] ^ d[187] ^ d[183] ^ d[182] ^ d[180] ^ d[179] ^ d[177] ^ d[175] ^ d[174] ^ d[169] ^ d[168] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[160] ^ d[159] ^ d[156] ^ d[155] ^ d[152] ^ d[150] ^ d[149] ^ d[148] ^ d[147] ^ d[146] ^ d[145] ^ d[144] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[136] ^ d[131] ^ d[127] ^ d[125] ^ d[122] ^ d[119] ^ d[117] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[108] ^ d[102] ^ d[100] ^ d[99] ^ d[92] ^ d[90] ^ d[88] ^ d[86] ^ d[85] ^ d[84] ^ d[81] ^ d[79] ^ d[78] ^ d[76] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[62] ^ d[60] ^ d[59] ^ d[56] ^ d[55] ^ d[53] ^ d[52] ^ d[46] ^ d[39] ^ d[37] ^ d[36] ^ d[32] ^ d[31] ^ d[30] ^ d[26] ^ d[24] ^ d[23] ^ d[16] ^ d[15] ^ d[12] ^ d[8] ^ d[4] ^ c[2] ^ c[7] ^ c[8] ^ c[10] ^ c[12] ^ c[13];
    newcrc[5] = d[1023] ^ d[1022] ^ d[1020] ^ d[1019] ^ d[1014] ^ d[1012] ^ d[1007] ^ d[1006] ^ d[1004] ^ d[1003] ^ d[1001] ^ d[1000] ^ d[999] ^ d[992] ^ d[990] ^ d[989] ^ d[987] ^ d[983] ^ d[982] ^ d[980] ^ d[976] ^ d[974] ^ d[973] ^ d[971] ^ d[970] ^ d[969] ^ d[967] ^ d[965] ^ d[964] ^ d[961] ^ d[956] ^ d[954] ^ d[952] ^ d[949] ^ d[948] ^ d[947] ^ d[945] ^ d[943] ^ d[940] ^ d[937] ^ d[929] ^ d[928] ^ d[927] ^ d[925] ^ d[923] ^ d[922] ^ d[921] ^ d[920] ^ d[918] ^ d[913] ^ d[912] ^ d[910] ^ d[904] ^ d[902] ^ d[901] ^ d[900] ^ d[899] ^ d[898] ^ d[895] ^ d[893] ^ d[892] ^ d[889] ^ d[888] ^ d[885] ^ d[883] ^ d[882] ^ d[881] ^ d[879] ^ d[878] ^ d[877] ^ d[876] ^ d[874] ^ d[873] ^ d[870] ^ d[869] ^ d[868] ^ d[865] ^ d[856] ^ d[854] ^ d[852] ^ d[851] ^ d[847] ^ d[846] ^ d[844] ^ d[841] ^ d[838] ^ d[834] ^ d[833] ^ d[832] ^ d[831] ^ d[830] ^ d[827] ^ d[822] ^ d[821] ^ d[820] ^ d[819] ^ d[815] ^ d[811] ^ d[809] ^ d[808] ^ d[807] ^ d[805] ^ d[803] ^ d[802] ^ d[800] ^ d[798] ^ d[796] ^ d[795] ^ d[793] ^ d[792] ^ d[791] ^ d[789] ^ d[786] ^ d[784] ^ d[783] ^ d[782] ^ d[779] ^ d[778] ^ d[777] ^ d[776] ^ d[775] ^ d[770] ^ d[768] ^ d[764] ^ d[763] ^ d[762] ^ d[761] ^ d[760] ^ d[757] ^ d[755] ^ d[754] ^ d[752] ^ d[751] ^ d[744] ^ d[743] ^ d[742] ^ d[741] ^ d[740] ^ d[739] ^ d[737] ^ d[734] ^ d[731] ^ d[730] ^ d[725] ^ d[724] ^ d[723] ^ d[722] ^ d[721] ^ d[720] ^ d[718] ^ d[717] ^ d[716] ^ d[714] ^ d[710] ^ d[709] ^ d[707] ^ d[705] ^ d[704] ^ d[702] ^ d[701] ^ d[699] ^ d[696] ^ d[695] ^ d[692] ^ d[688] ^ d[686] ^ d[685] ^ d[684] ^ d[683] ^ d[681] ^ d[680] ^ d[678] ^ d[676] ^ d[675] ^ d[674] ^ d[669] ^ d[667] ^ d[666] ^ d[665] ^ d[664] ^ d[663] ^ d[662] ^ d[661] ^ d[656] ^ d[655] ^ d[654] ^ d[652] ^ d[651] ^ d[650] ^ d[649] ^ d[648] ^ d[642] ^ d[635] ^ d[634] ^ d[633] ^ d[632] ^ d[629] ^ d[628] ^ d[627] ^ d[626] ^ d[624] ^ d[620] ^ d[618] ^ d[614] ^ d[611] ^ d[610] ^ d[609] ^ d[605] ^ d[600] ^ d[599] ^ d[597] ^ d[592] ^ d[589] ^ d[588] ^ d[585] ^ d[581] ^ d[577] ^ d[576] ^ d[571] ^ d[566] ^ d[564] ^ d[560] ^ d[554] ^ d[552] ^ d[550] ^ d[549] ^ d[547] ^ d[545] ^ d[537] ^ d[536] ^ d[535] ^ d[534] ^ d[532] ^ d[530] ^ d[527] ^ d[524] ^ d[523] ^ d[521] ^ d[518] ^ d[515] ^ d[514] ^ d[513] ^ d[512] ^ d[510] ^ d[506] ^ d[503] ^ d[500] ^ d[499] ^ d[498] ^ d[497] ^ d[496] ^ d[495] ^ d[494] ^ d[493] ^ d[492] ^ d[489] ^ d[487] ^ d[486] ^ d[485] ^ d[484] ^ d[482] ^ d[481] ^ d[480] ^ d[478] ^ d[477] ^ d[474] ^ d[473] ^ d[471] ^ d[469] ^ d[468] ^ d[466] ^ d[463] ^ d[461] ^ d[459] ^ d[455] ^ d[453] ^ d[452] ^ d[451] ^ d[449] ^ d[448] ^ d[447] ^ d[446] ^ d[445] ^ d[444] ^ d[443] ^ d[442] ^ d[439] ^ d[438] ^ d[437] ^ d[433] ^ d[432] ^ d[429] ^ d[427] ^ d[425] ^ d[424] ^ d[423] ^ d[419] ^ d[418] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[411] ^ d[410] ^ d[407] ^ d[405] ^ d[404] ^ d[402] ^ d[401] ^ d[400] ^ d[399] ^ d[395] ^ d[393] ^ d[392] ^ d[391] ^ d[388] ^ d[385] ^ d[384] ^ d[383] ^ d[381] ^ d[379] ^ d[378] ^ d[377] ^ d[376] ^ d[375] ^ d[374] ^ d[372] ^ d[370] ^ d[369] ^ d[368] ^ d[367] ^ d[366] ^ d[365] ^ d[363] ^ d[362] ^ d[360] ^ d[359] ^ d[358] ^ d[354] ^ d[353] ^ d[352] ^ d[347] ^ d[344] ^ d[343] ^ d[342] ^ d[341] ^ d[340] ^ d[339] ^ d[334] ^ d[332] ^ d[330] ^ d[327] ^ d[326] ^ d[324] ^ d[323] ^ d[321] ^ d[320] ^ d[319] ^ d[318] ^ d[314] ^ d[313] ^ d[312] ^ d[310] ^ d[308] ^ d[307] ^ d[306] ^ d[304] ^ d[302] ^ d[300] ^ d[299] ^ d[294] ^ d[291] ^ d[289] ^ d[287] ^ d[283] ^ d[279] ^ d[277] ^ d[274] ^ d[273] ^ d[272] ^ d[269] ^ d[268] ^ d[267] ^ d[265] ^ d[264] ^ d[259] ^ d[258] ^ d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[247] ^ d[245] ^ d[242] ^ d[241] ^ d[240] ^ d[236] ^ d[235] ^ d[234] ^ d[233] ^ d[229] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[217] ^ d[214] ^ d[211] ^ d[208] ^ d[207] ^ d[205] ^ d[203] ^ d[201] ^ d[200] ^ d[199] ^ d[195] ^ d[194] ^ d[193] ^ d[192] ^ d[190] ^ d[189] ^ d[187] ^ d[181] ^ d[180] ^ d[179] ^ d[173] ^ d[171] ^ d[169] ^ d[167] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[160] ^ d[159] ^ d[158] ^ d[157] ^ d[155] ^ d[153] ^ d[152] ^ d[150] ^ d[149] ^ d[147] ^ d[140] ^ d[139] ^ d[138] ^ d[136] ^ d[128] ^ d[127] ^ d[126] ^ d[121] ^ d[120] ^ d[114] ^ d[112] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[101] ^ d[100] ^ d[98] ^ d[96] ^ d[95] ^ d[93] ^ d[91] ^ d[89] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[81] ^ d[79] ^ d[74] ^ d[71] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[64] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[42] ^ d[40] ^ d[38] ^ d[37] ^ d[35] ^ d[31] ^ d[28] ^ d[26] ^ d[25] ^ d[24] ^ d[22] ^ d[20] ^ d[19] ^ d[17] ^ d[16] ^ d[13] ^ d[12] ^ d[11] ^ d[9] ^ d[8] ^ d[5] ^ d[4] ^ d[0] ^ c[4] ^ c[6] ^ c[11] ^ c[12] ^ c[14] ^ c[15];
    newcrc[6] = d[1023] ^ d[1021] ^ d[1020] ^ d[1015] ^ d[1013] ^ d[1008] ^ d[1007] ^ d[1005] ^ d[1004] ^ d[1002] ^ d[1001] ^ d[1000] ^ d[993] ^ d[991] ^ d[990] ^ d[988] ^ d[984] ^ d[983] ^ d[981] ^ d[977] ^ d[975] ^ d[974] ^ d[972] ^ d[971] ^ d[970] ^ d[968] ^ d[966] ^ d[965] ^ d[962] ^ d[957] ^ d[955] ^ d[953] ^ d[950] ^ d[949] ^ d[948] ^ d[946] ^ d[944] ^ d[941] ^ d[938] ^ d[930] ^ d[929] ^ d[928] ^ d[926] ^ d[924] ^ d[923] ^ d[922] ^ d[921] ^ d[919] ^ d[914] ^ d[913] ^ d[911] ^ d[905] ^ d[903] ^ d[902] ^ d[901] ^ d[900] ^ d[899] ^ d[896] ^ d[894] ^ d[893] ^ d[890] ^ d[889] ^ d[886] ^ d[884] ^ d[883] ^ d[882] ^ d[880] ^ d[879] ^ d[878] ^ d[877] ^ d[875] ^ d[874] ^ d[871] ^ d[870] ^ d[869] ^ d[866] ^ d[857] ^ d[855] ^ d[853] ^ d[852] ^ d[848] ^ d[847] ^ d[845] ^ d[842] ^ d[839] ^ d[835] ^ d[834] ^ d[833] ^ d[832] ^ d[831] ^ d[828] ^ d[823] ^ d[822] ^ d[821] ^ d[820] ^ d[816] ^ d[812] ^ d[810] ^ d[809] ^ d[808] ^ d[806] ^ d[804] ^ d[803] ^ d[801] ^ d[799] ^ d[797] ^ d[796] ^ d[794] ^ d[793] ^ d[792] ^ d[790] ^ d[787] ^ d[785] ^ d[784] ^ d[783] ^ d[780] ^ d[779] ^ d[778] ^ d[777] ^ d[776] ^ d[771] ^ d[769] ^ d[765] ^ d[764] ^ d[763] ^ d[762] ^ d[761] ^ d[758] ^ d[756] ^ d[755] ^ d[753] ^ d[752] ^ d[745] ^ d[744] ^ d[743] ^ d[742] ^ d[741] ^ d[740] ^ d[738] ^ d[735] ^ d[732] ^ d[731] ^ d[726] ^ d[725] ^ d[724] ^ d[723] ^ d[722] ^ d[721] ^ d[719] ^ d[718] ^ d[717] ^ d[715] ^ d[711] ^ d[710] ^ d[708] ^ d[706] ^ d[705] ^ d[703] ^ d[702] ^ d[700] ^ d[697] ^ d[696] ^ d[693] ^ d[689] ^ d[687] ^ d[686] ^ d[685] ^ d[684] ^ d[682] ^ d[681] ^ d[679] ^ d[677] ^ d[676] ^ d[675] ^ d[670] ^ d[668] ^ d[667] ^ d[666] ^ d[665] ^ d[664] ^ d[663] ^ d[662] ^ d[657] ^ d[656] ^ d[655] ^ d[653] ^ d[652] ^ d[651] ^ d[650] ^ d[649] ^ d[643] ^ d[636] ^ d[635] ^ d[634] ^ d[633] ^ d[630] ^ d[629] ^ d[628] ^ d[627] ^ d[625] ^ d[621] ^ d[619] ^ d[615] ^ d[612] ^ d[611] ^ d[610] ^ d[606] ^ d[601] ^ d[600] ^ d[598] ^ d[593] ^ d[590] ^ d[589] ^ d[586] ^ d[582] ^ d[578] ^ d[577] ^ d[572] ^ d[567] ^ d[565] ^ d[561] ^ d[555] ^ d[553] ^ d[551] ^ d[550] ^ d[548] ^ d[546] ^ d[538] ^ d[537] ^ d[536] ^ d[535] ^ d[533] ^ d[531] ^ d[528] ^ d[525] ^ d[524] ^ d[522] ^ d[519] ^ d[516] ^ d[515] ^ d[514] ^ d[513] ^ d[511] ^ d[507] ^ d[504] ^ d[501] ^ d[500] ^ d[499] ^ d[498] ^ d[497] ^ d[496] ^ d[495] ^ d[494] ^ d[493] ^ d[490] ^ d[488] ^ d[487] ^ d[486] ^ d[485] ^ d[483] ^ d[482] ^ d[481] ^ d[479] ^ d[478] ^ d[475] ^ d[474] ^ d[472] ^ d[470] ^ d[469] ^ d[467] ^ d[464] ^ d[462] ^ d[460] ^ d[456] ^ d[454] ^ d[453] ^ d[452] ^ d[450] ^ d[449] ^ d[448] ^ d[447] ^ d[446] ^ d[445] ^ d[444] ^ d[443] ^ d[440] ^ d[439] ^ d[438] ^ d[434] ^ d[433] ^ d[430] ^ d[428] ^ d[426] ^ d[425] ^ d[424] ^ d[420] ^ d[419] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[411] ^ d[408] ^ d[406] ^ d[405] ^ d[403] ^ d[402] ^ d[401] ^ d[400] ^ d[396] ^ d[394] ^ d[393] ^ d[392] ^ d[389] ^ d[386] ^ d[385] ^ d[384] ^ d[382] ^ d[380] ^ d[379] ^ d[378] ^ d[377] ^ d[376] ^ d[375] ^ d[373] ^ d[371] ^ d[370] ^ d[369] ^ d[368] ^ d[367] ^ d[366] ^ d[364] ^ d[363] ^ d[361] ^ d[360] ^ d[359] ^ d[355] ^ d[354] ^ d[353] ^ d[348] ^ d[345] ^ d[344] ^ d[343] ^ d[342] ^ d[341] ^ d[340] ^ d[335] ^ d[333] ^ d[331] ^ d[328] ^ d[327] ^ d[325] ^ d[324] ^ d[322] ^ d[321] ^ d[320] ^ d[319] ^ d[315] ^ d[314] ^ d[313] ^ d[311] ^ d[309] ^ d[308] ^ d[307] ^ d[305] ^ d[303] ^ d[301] ^ d[300] ^ d[295] ^ d[292] ^ d[290] ^ d[288] ^ d[284] ^ d[280] ^ d[278] ^ d[275] ^ d[274] ^ d[273] ^ d[270] ^ d[269] ^ d[268] ^ d[266] ^ d[265] ^ d[260] ^ d[259] ^ d[256] ^ d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[248] ^ d[246] ^ d[243] ^ d[242] ^ d[241] ^ d[237] ^ d[236] ^ d[235] ^ d[234] ^ d[230] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[218] ^ d[215] ^ d[212] ^ d[209] ^ d[208] ^ d[206] ^ d[204] ^ d[202] ^ d[201] ^ d[200] ^ d[196] ^ d[195] ^ d[194] ^ d[193] ^ d[191] ^ d[190] ^ d[188] ^ d[182] ^ d[181] ^ d[180] ^ d[174] ^ d[172] ^ d[170] ^ d[168] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[161] ^ d[160] ^ d[159] ^ d[158] ^ d[156] ^ d[154] ^ d[153] ^ d[151] ^ d[150] ^ d[148] ^ d[141] ^ d[140] ^ d[139] ^ d[137] ^ d[129] ^ d[128] ^ d[127] ^ d[122] ^ d[121] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[99] ^ d[97] ^ d[96] ^ d[94] ^ d[92] ^ d[90] ^ d[89] ^ d[88] ^ d[86] ^ d[85] ^ d[82] ^ d[80] ^ d[75] ^ d[72] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[62] ^ d[61] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[50] ^ d[49] ^ d[48] ^ d[43] ^ d[41] ^ d[39] ^ d[38] ^ d[36] ^ d[32] ^ d[29] ^ d[27] ^ d[26] ^ d[25] ^ d[23] ^ d[21] ^ d[20] ^ d[18] ^ d[17] ^ d[14] ^ d[13] ^ d[12] ^ d[10] ^ d[9] ^ d[6] ^ d[5] ^ d[1] ^ c[0] ^ c[5] ^ c[7] ^ c[12] ^ c[13] ^ c[15];
    newcrc[7] = d[1022] ^ d[1021] ^ d[1016] ^ d[1014] ^ d[1009] ^ d[1008] ^ d[1006] ^ d[1005] ^ d[1003] ^ d[1002] ^ d[1001] ^ d[994] ^ d[992] ^ d[991] ^ d[989] ^ d[985] ^ d[984] ^ d[982] ^ d[978] ^ d[976] ^ d[975] ^ d[973] ^ d[972] ^ d[971] ^ d[969] ^ d[967] ^ d[966] ^ d[963] ^ d[958] ^ d[956] ^ d[954] ^ d[951] ^ d[950] ^ d[949] ^ d[947] ^ d[945] ^ d[942] ^ d[939] ^ d[931] ^ d[930] ^ d[929] ^ d[927] ^ d[925] ^ d[924] ^ d[923] ^ d[922] ^ d[920] ^ d[915] ^ d[914] ^ d[912] ^ d[906] ^ d[904] ^ d[903] ^ d[902] ^ d[901] ^ d[900] ^ d[897] ^ d[895] ^ d[894] ^ d[891] ^ d[890] ^ d[887] ^ d[885] ^ d[884] ^ d[883] ^ d[881] ^ d[880] ^ d[879] ^ d[878] ^ d[876] ^ d[875] ^ d[872] ^ d[871] ^ d[870] ^ d[867] ^ d[858] ^ d[856] ^ d[854] ^ d[853] ^ d[849] ^ d[848] ^ d[846] ^ d[843] ^ d[840] ^ d[836] ^ d[835] ^ d[834] ^ d[833] ^ d[832] ^ d[829] ^ d[824] ^ d[823] ^ d[822] ^ d[821] ^ d[817] ^ d[813] ^ d[811] ^ d[810] ^ d[809] ^ d[807] ^ d[805] ^ d[804] ^ d[802] ^ d[800] ^ d[798] ^ d[797] ^ d[795] ^ d[794] ^ d[793] ^ d[791] ^ d[788] ^ d[786] ^ d[785] ^ d[784] ^ d[781] ^ d[780] ^ d[779] ^ d[778] ^ d[777] ^ d[772] ^ d[770] ^ d[766] ^ d[765] ^ d[764] ^ d[763] ^ d[762] ^ d[759] ^ d[757] ^ d[756] ^ d[754] ^ d[753] ^ d[746] ^ d[745] ^ d[744] ^ d[743] ^ d[742] ^ d[741] ^ d[739] ^ d[736] ^ d[733] ^ d[732] ^ d[727] ^ d[726] ^ d[725] ^ d[724] ^ d[723] ^ d[722] ^ d[720] ^ d[719] ^ d[718] ^ d[716] ^ d[712] ^ d[711] ^ d[709] ^ d[707] ^ d[706] ^ d[704] ^ d[703] ^ d[701] ^ d[698] ^ d[697] ^ d[694] ^ d[690] ^ d[688] ^ d[687] ^ d[686] ^ d[685] ^ d[683] ^ d[682] ^ d[680] ^ d[678] ^ d[677] ^ d[676] ^ d[671] ^ d[669] ^ d[668] ^ d[667] ^ d[666] ^ d[665] ^ d[664] ^ d[663] ^ d[658] ^ d[657] ^ d[656] ^ d[654] ^ d[653] ^ d[652] ^ d[651] ^ d[650] ^ d[644] ^ d[637] ^ d[636] ^ d[635] ^ d[634] ^ d[631] ^ d[630] ^ d[629] ^ d[628] ^ d[626] ^ d[622] ^ d[620] ^ d[616] ^ d[613] ^ d[612] ^ d[611] ^ d[607] ^ d[602] ^ d[601] ^ d[599] ^ d[594] ^ d[591] ^ d[590] ^ d[587] ^ d[583] ^ d[579] ^ d[578] ^ d[573] ^ d[568] ^ d[566] ^ d[562] ^ d[556] ^ d[554] ^ d[552] ^ d[551] ^ d[549] ^ d[547] ^ d[539] ^ d[538] ^ d[537] ^ d[536] ^ d[534] ^ d[532] ^ d[529] ^ d[526] ^ d[525] ^ d[523] ^ d[520] ^ d[517] ^ d[516] ^ d[515] ^ d[514] ^ d[512] ^ d[508] ^ d[505] ^ d[502] ^ d[501] ^ d[500] ^ d[499] ^ d[498] ^ d[497] ^ d[496] ^ d[495] ^ d[494] ^ d[491] ^ d[489] ^ d[488] ^ d[487] ^ d[486] ^ d[484] ^ d[483] ^ d[482] ^ d[480] ^ d[479] ^ d[476] ^ d[475] ^ d[473] ^ d[471] ^ d[470] ^ d[468] ^ d[465] ^ d[463] ^ d[461] ^ d[457] ^ d[455] ^ d[454] ^ d[453] ^ d[451] ^ d[450] ^ d[449] ^ d[448] ^ d[447] ^ d[446] ^ d[445] ^ d[444] ^ d[441] ^ d[440] ^ d[439] ^ d[435] ^ d[434] ^ d[431] ^ d[429] ^ d[427] ^ d[426] ^ d[425] ^ d[421] ^ d[420] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[412] ^ d[409] ^ d[407] ^ d[406] ^ d[404] ^ d[403] ^ d[402] ^ d[401] ^ d[397] ^ d[395] ^ d[394] ^ d[393] ^ d[390] ^ d[387] ^ d[386] ^ d[385] ^ d[383] ^ d[381] ^ d[380] ^ d[379] ^ d[378] ^ d[377] ^ d[376] ^ d[374] ^ d[372] ^ d[371] ^ d[370] ^ d[369] ^ d[368] ^ d[367] ^ d[365] ^ d[364] ^ d[362] ^ d[361] ^ d[360] ^ d[356] ^ d[355] ^ d[354] ^ d[349] ^ d[346] ^ d[345] ^ d[344] ^ d[343] ^ d[342] ^ d[341] ^ d[336] ^ d[334] ^ d[332] ^ d[329] ^ d[328] ^ d[326] ^ d[325] ^ d[323] ^ d[322] ^ d[321] ^ d[320] ^ d[316] ^ d[315] ^ d[314] ^ d[312] ^ d[310] ^ d[309] ^ d[308] ^ d[306] ^ d[304] ^ d[302] ^ d[301] ^ d[296] ^ d[293] ^ d[291] ^ d[289] ^ d[285] ^ d[281] ^ d[279] ^ d[276] ^ d[275] ^ d[274] ^ d[271] ^ d[270] ^ d[269] ^ d[267] ^ d[266] ^ d[261] ^ d[260] ^ d[257] ^ d[256] ^ d[255] ^ d[253] ^ d[252] ^ d[249] ^ d[247] ^ d[244] ^ d[243] ^ d[242] ^ d[238] ^ d[237] ^ d[236] ^ d[235] ^ d[231] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[219] ^ d[216] ^ d[213] ^ d[210] ^ d[209] ^ d[207] ^ d[205] ^ d[203] ^ d[202] ^ d[201] ^ d[197] ^ d[196] ^ d[195] ^ d[194] ^ d[192] ^ d[191] ^ d[189] ^ d[183] ^ d[182] ^ d[181] ^ d[175] ^ d[173] ^ d[171] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[164] ^ d[162] ^ d[161] ^ d[160] ^ d[159] ^ d[157] ^ d[155] ^ d[154] ^ d[152] ^ d[151] ^ d[149] ^ d[142] ^ d[141] ^ d[140] ^ d[138] ^ d[130] ^ d[129] ^ d[128] ^ d[123] ^ d[122] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[100] ^ d[98] ^ d[97] ^ d[95] ^ d[93] ^ d[91] ^ d[90] ^ d[89] ^ d[87] ^ d[86] ^ d[83] ^ d[81] ^ d[76] ^ d[73] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[44] ^ d[42] ^ d[40] ^ d[39] ^ d[37] ^ d[33] ^ d[30] ^ d[28] ^ d[27] ^ d[26] ^ d[24] ^ d[22] ^ d[21] ^ d[19] ^ d[18] ^ d[15] ^ d[14] ^ d[13] ^ d[11] ^ d[10] ^ d[7] ^ d[6] ^ d[2] ^ c[0] ^ c[1] ^ c[6] ^ c[8] ^ c[13] ^ c[14];
    newcrc[8] = d[1023] ^ d[1022] ^ d[1017] ^ d[1015] ^ d[1010] ^ d[1009] ^ d[1007] ^ d[1006] ^ d[1004] ^ d[1003] ^ d[1002] ^ d[995] ^ d[993] ^ d[992] ^ d[990] ^ d[986] ^ d[985] ^ d[983] ^ d[979] ^ d[977] ^ d[976] ^ d[974] ^ d[973] ^ d[972] ^ d[970] ^ d[968] ^ d[967] ^ d[964] ^ d[959] ^ d[957] ^ d[955] ^ d[952] ^ d[951] ^ d[950] ^ d[948] ^ d[946] ^ d[943] ^ d[940] ^ d[932] ^ d[931] ^ d[930] ^ d[928] ^ d[926] ^ d[925] ^ d[924] ^ d[923] ^ d[921] ^ d[916] ^ d[915] ^ d[913] ^ d[907] ^ d[905] ^ d[904] ^ d[903] ^ d[902] ^ d[901] ^ d[898] ^ d[896] ^ d[895] ^ d[892] ^ d[891] ^ d[888] ^ d[886] ^ d[885] ^ d[884] ^ d[882] ^ d[881] ^ d[880] ^ d[879] ^ d[877] ^ d[876] ^ d[873] ^ d[872] ^ d[871] ^ d[868] ^ d[859] ^ d[857] ^ d[855] ^ d[854] ^ d[850] ^ d[849] ^ d[847] ^ d[844] ^ d[841] ^ d[837] ^ d[836] ^ d[835] ^ d[834] ^ d[833] ^ d[830] ^ d[825] ^ d[824] ^ d[823] ^ d[822] ^ d[818] ^ d[814] ^ d[812] ^ d[811] ^ d[810] ^ d[808] ^ d[806] ^ d[805] ^ d[803] ^ d[801] ^ d[799] ^ d[798] ^ d[796] ^ d[795] ^ d[794] ^ d[792] ^ d[789] ^ d[787] ^ d[786] ^ d[785] ^ d[782] ^ d[781] ^ d[780] ^ d[779] ^ d[778] ^ d[773] ^ d[771] ^ d[767] ^ d[766] ^ d[765] ^ d[764] ^ d[763] ^ d[760] ^ d[758] ^ d[757] ^ d[755] ^ d[754] ^ d[747] ^ d[746] ^ d[745] ^ d[744] ^ d[743] ^ d[742] ^ d[740] ^ d[737] ^ d[734] ^ d[733] ^ d[728] ^ d[727] ^ d[726] ^ d[725] ^ d[724] ^ d[723] ^ d[721] ^ d[720] ^ d[719] ^ d[717] ^ d[713] ^ d[712] ^ d[710] ^ d[708] ^ d[707] ^ d[705] ^ d[704] ^ d[702] ^ d[699] ^ d[698] ^ d[695] ^ d[691] ^ d[689] ^ d[688] ^ d[687] ^ d[686] ^ d[684] ^ d[683] ^ d[681] ^ d[679] ^ d[678] ^ d[677] ^ d[672] ^ d[670] ^ d[669] ^ d[668] ^ d[667] ^ d[666] ^ d[665] ^ d[664] ^ d[659] ^ d[658] ^ d[657] ^ d[655] ^ d[654] ^ d[653] ^ d[652] ^ d[651] ^ d[645] ^ d[638] ^ d[637] ^ d[636] ^ d[635] ^ d[632] ^ d[631] ^ d[630] ^ d[629] ^ d[627] ^ d[623] ^ d[621] ^ d[617] ^ d[614] ^ d[613] ^ d[612] ^ d[608] ^ d[603] ^ d[602] ^ d[600] ^ d[595] ^ d[592] ^ d[591] ^ d[588] ^ d[584] ^ d[580] ^ d[579] ^ d[574] ^ d[569] ^ d[567] ^ d[563] ^ d[557] ^ d[555] ^ d[553] ^ d[552] ^ d[550] ^ d[548] ^ d[540] ^ d[539] ^ d[538] ^ d[537] ^ d[535] ^ d[533] ^ d[530] ^ d[527] ^ d[526] ^ d[524] ^ d[521] ^ d[518] ^ d[517] ^ d[516] ^ d[515] ^ d[513] ^ d[509] ^ d[506] ^ d[503] ^ d[502] ^ d[501] ^ d[500] ^ d[499] ^ d[498] ^ d[497] ^ d[496] ^ d[495] ^ d[492] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[485] ^ d[484] ^ d[483] ^ d[481] ^ d[480] ^ d[477] ^ d[476] ^ d[474] ^ d[472] ^ d[471] ^ d[469] ^ d[466] ^ d[464] ^ d[462] ^ d[458] ^ d[456] ^ d[455] ^ d[454] ^ d[452] ^ d[451] ^ d[450] ^ d[449] ^ d[448] ^ d[447] ^ d[446] ^ d[445] ^ d[442] ^ d[441] ^ d[440] ^ d[436] ^ d[435] ^ d[432] ^ d[430] ^ d[428] ^ d[427] ^ d[426] ^ d[422] ^ d[421] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[413] ^ d[410] ^ d[408] ^ d[407] ^ d[405] ^ d[404] ^ d[403] ^ d[402] ^ d[398] ^ d[396] ^ d[395] ^ d[394] ^ d[391] ^ d[388] ^ d[387] ^ d[386] ^ d[384] ^ d[382] ^ d[381] ^ d[380] ^ d[379] ^ d[378] ^ d[377] ^ d[375] ^ d[373] ^ d[372] ^ d[371] ^ d[370] ^ d[369] ^ d[368] ^ d[366] ^ d[365] ^ d[363] ^ d[362] ^ d[361] ^ d[357] ^ d[356] ^ d[355] ^ d[350] ^ d[347] ^ d[346] ^ d[345] ^ d[344] ^ d[343] ^ d[342] ^ d[337] ^ d[335] ^ d[333] ^ d[330] ^ d[329] ^ d[327] ^ d[326] ^ d[324] ^ d[323] ^ d[322] ^ d[321] ^ d[317] ^ d[316] ^ d[315] ^ d[313] ^ d[311] ^ d[310] ^ d[309] ^ d[307] ^ d[305] ^ d[303] ^ d[302] ^ d[297] ^ d[294] ^ d[292] ^ d[290] ^ d[286] ^ d[282] ^ d[280] ^ d[277] ^ d[276] ^ d[275] ^ d[272] ^ d[271] ^ d[270] ^ d[268] ^ d[267] ^ d[262] ^ d[261] ^ d[258] ^ d[257] ^ d[256] ^ d[254] ^ d[253] ^ d[250] ^ d[248] ^ d[245] ^ d[244] ^ d[243] ^ d[239] ^ d[238] ^ d[237] ^ d[236] ^ d[232] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[220] ^ d[217] ^ d[214] ^ d[211] ^ d[210] ^ d[208] ^ d[206] ^ d[204] ^ d[203] ^ d[202] ^ d[198] ^ d[197] ^ d[196] ^ d[195] ^ d[193] ^ d[192] ^ d[190] ^ d[184] ^ d[183] ^ d[182] ^ d[176] ^ d[174] ^ d[172] ^ d[170] ^ d[169] ^ d[168] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[161] ^ d[160] ^ d[158] ^ d[156] ^ d[155] ^ d[153] ^ d[152] ^ d[150] ^ d[143] ^ d[142] ^ d[141] ^ d[139] ^ d[131] ^ d[130] ^ d[129] ^ d[124] ^ d[123] ^ d[117] ^ d[115] ^ d[114] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[94] ^ d[92] ^ d[91] ^ d[90] ^ d[88] ^ d[87] ^ d[84] ^ d[82] ^ d[77] ^ d[74] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[64] ^ d[63] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[45] ^ d[43] ^ d[41] ^ d[40] ^ d[38] ^ d[34] ^ d[31] ^ d[29] ^ d[28] ^ d[27] ^ d[25] ^ d[23] ^ d[22] ^ d[20] ^ d[19] ^ d[16] ^ d[15] ^ d[14] ^ d[12] ^ d[11] ^ d[8] ^ d[7] ^ d[3] ^ c[1] ^ c[2] ^ c[7] ^ c[9] ^ c[14] ^ c[15];
    newcrc[9] = d[1023] ^ d[1018] ^ d[1016] ^ d[1011] ^ d[1010] ^ d[1008] ^ d[1007] ^ d[1005] ^ d[1004] ^ d[1003] ^ d[996] ^ d[994] ^ d[993] ^ d[991] ^ d[987] ^ d[986] ^ d[984] ^ d[980] ^ d[978] ^ d[977] ^ d[975] ^ d[974] ^ d[973] ^ d[971] ^ d[969] ^ d[968] ^ d[965] ^ d[960] ^ d[958] ^ d[956] ^ d[953] ^ d[952] ^ d[951] ^ d[949] ^ d[947] ^ d[944] ^ d[941] ^ d[933] ^ d[932] ^ d[931] ^ d[929] ^ d[927] ^ d[926] ^ d[925] ^ d[924] ^ d[922] ^ d[917] ^ d[916] ^ d[914] ^ d[908] ^ d[906] ^ d[905] ^ d[904] ^ d[903] ^ d[902] ^ d[899] ^ d[897] ^ d[896] ^ d[893] ^ d[892] ^ d[889] ^ d[887] ^ d[886] ^ d[885] ^ d[883] ^ d[882] ^ d[881] ^ d[880] ^ d[878] ^ d[877] ^ d[874] ^ d[873] ^ d[872] ^ d[869] ^ d[860] ^ d[858] ^ d[856] ^ d[855] ^ d[851] ^ d[850] ^ d[848] ^ d[845] ^ d[842] ^ d[838] ^ d[837] ^ d[836] ^ d[835] ^ d[834] ^ d[831] ^ d[826] ^ d[825] ^ d[824] ^ d[823] ^ d[819] ^ d[815] ^ d[813] ^ d[812] ^ d[811] ^ d[809] ^ d[807] ^ d[806] ^ d[804] ^ d[802] ^ d[800] ^ d[799] ^ d[797] ^ d[796] ^ d[795] ^ d[793] ^ d[790] ^ d[788] ^ d[787] ^ d[786] ^ d[783] ^ d[782] ^ d[781] ^ d[780] ^ d[779] ^ d[774] ^ d[772] ^ d[768] ^ d[767] ^ d[766] ^ d[765] ^ d[764] ^ d[761] ^ d[759] ^ d[758] ^ d[756] ^ d[755] ^ d[748] ^ d[747] ^ d[746] ^ d[745] ^ d[744] ^ d[743] ^ d[741] ^ d[738] ^ d[735] ^ d[734] ^ d[729] ^ d[728] ^ d[727] ^ d[726] ^ d[725] ^ d[724] ^ d[722] ^ d[721] ^ d[720] ^ d[718] ^ d[714] ^ d[713] ^ d[711] ^ d[709] ^ d[708] ^ d[706] ^ d[705] ^ d[703] ^ d[700] ^ d[699] ^ d[696] ^ d[692] ^ d[690] ^ d[689] ^ d[688] ^ d[687] ^ d[685] ^ d[684] ^ d[682] ^ d[680] ^ d[679] ^ d[678] ^ d[673] ^ d[671] ^ d[670] ^ d[669] ^ d[668] ^ d[667] ^ d[666] ^ d[665] ^ d[660] ^ d[659] ^ d[658] ^ d[656] ^ d[655] ^ d[654] ^ d[653] ^ d[652] ^ d[646] ^ d[639] ^ d[638] ^ d[637] ^ d[636] ^ d[633] ^ d[632] ^ d[631] ^ d[630] ^ d[628] ^ d[624] ^ d[622] ^ d[618] ^ d[615] ^ d[614] ^ d[613] ^ d[609] ^ d[604] ^ d[603] ^ d[601] ^ d[596] ^ d[593] ^ d[592] ^ d[589] ^ d[585] ^ d[581] ^ d[580] ^ d[575] ^ d[570] ^ d[568] ^ d[564] ^ d[558] ^ d[556] ^ d[554] ^ d[553] ^ d[551] ^ d[549] ^ d[541] ^ d[540] ^ d[539] ^ d[538] ^ d[536] ^ d[534] ^ d[531] ^ d[528] ^ d[527] ^ d[525] ^ d[522] ^ d[519] ^ d[518] ^ d[517] ^ d[516] ^ d[514] ^ d[510] ^ d[507] ^ d[504] ^ d[503] ^ d[502] ^ d[501] ^ d[500] ^ d[499] ^ d[498] ^ d[497] ^ d[496] ^ d[493] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[486] ^ d[485] ^ d[484] ^ d[482] ^ d[481] ^ d[478] ^ d[477] ^ d[475] ^ d[473] ^ d[472] ^ d[470] ^ d[467] ^ d[465] ^ d[463] ^ d[459] ^ d[457] ^ d[456] ^ d[455] ^ d[453] ^ d[452] ^ d[451] ^ d[450] ^ d[449] ^ d[448] ^ d[447] ^ d[446] ^ d[443] ^ d[442] ^ d[441] ^ d[437] ^ d[436] ^ d[433] ^ d[431] ^ d[429] ^ d[428] ^ d[427] ^ d[423] ^ d[422] ^ d[420] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[414] ^ d[411] ^ d[409] ^ d[408] ^ d[406] ^ d[405] ^ d[404] ^ d[403] ^ d[399] ^ d[397] ^ d[396] ^ d[395] ^ d[392] ^ d[389] ^ d[388] ^ d[387] ^ d[385] ^ d[383] ^ d[382] ^ d[381] ^ d[380] ^ d[379] ^ d[378] ^ d[376] ^ d[374] ^ d[373] ^ d[372] ^ d[371] ^ d[370] ^ d[369] ^ d[367] ^ d[366] ^ d[364] ^ d[363] ^ d[362] ^ d[358] ^ d[357] ^ d[356] ^ d[351] ^ d[348] ^ d[347] ^ d[346] ^ d[345] ^ d[344] ^ d[343] ^ d[338] ^ d[336] ^ d[334] ^ d[331] ^ d[330] ^ d[328] ^ d[327] ^ d[325] ^ d[324] ^ d[323] ^ d[322] ^ d[318] ^ d[317] ^ d[316] ^ d[314] ^ d[312] ^ d[311] ^ d[310] ^ d[308] ^ d[306] ^ d[304] ^ d[303] ^ d[298] ^ d[295] ^ d[293] ^ d[291] ^ d[287] ^ d[283] ^ d[281] ^ d[278] ^ d[277] ^ d[276] ^ d[273] ^ d[272] ^ d[271] ^ d[269] ^ d[268] ^ d[263] ^ d[262] ^ d[259] ^ d[258] ^ d[257] ^ d[255] ^ d[254] ^ d[251] ^ d[249] ^ d[246] ^ d[245] ^ d[244] ^ d[240] ^ d[239] ^ d[238] ^ d[237] ^ d[233] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[221] ^ d[218] ^ d[215] ^ d[212] ^ d[211] ^ d[209] ^ d[207] ^ d[205] ^ d[204] ^ d[203] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[194] ^ d[193] ^ d[191] ^ d[185] ^ d[184] ^ d[183] ^ d[177] ^ d[175] ^ d[173] ^ d[171] ^ d[170] ^ d[169] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[159] ^ d[157] ^ d[156] ^ d[154] ^ d[153] ^ d[151] ^ d[144] ^ d[143] ^ d[142] ^ d[140] ^ d[132] ^ d[131] ^ d[130] ^ d[125] ^ d[124] ^ d[118] ^ d[116] ^ d[115] ^ d[114] ^ d[112] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[102] ^ d[100] ^ d[99] ^ d[97] ^ d[95] ^ d[93] ^ d[92] ^ d[91] ^ d[89] ^ d[88] ^ d[85] ^ d[83] ^ d[78] ^ d[75] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[65] ^ d[64] ^ d[62] ^ d[61] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[46] ^ d[44] ^ d[42] ^ d[41] ^ d[39] ^ d[35] ^ d[32] ^ d[30] ^ d[29] ^ d[28] ^ d[26] ^ d[24] ^ d[23] ^ d[21] ^ d[20] ^ d[17] ^ d[16] ^ d[15] ^ d[13] ^ d[12] ^ d[9] ^ d[8] ^ d[4] ^ c[0] ^ c[2] ^ c[3] ^ c[8] ^ c[10] ^ c[15];
    newcrc[10] = d[1019] ^ d[1017] ^ d[1012] ^ d[1011] ^ d[1009] ^ d[1008] ^ d[1006] ^ d[1005] ^ d[1004] ^ d[997] ^ d[995] ^ d[994] ^ d[992] ^ d[988] ^ d[987] ^ d[985] ^ d[981] ^ d[979] ^ d[978] ^ d[976] ^ d[975] ^ d[974] ^ d[972] ^ d[970] ^ d[969] ^ d[966] ^ d[961] ^ d[959] ^ d[957] ^ d[954] ^ d[953] ^ d[952] ^ d[950] ^ d[948] ^ d[945] ^ d[942] ^ d[934] ^ d[933] ^ d[932] ^ d[930] ^ d[928] ^ d[927] ^ d[926] ^ d[925] ^ d[923] ^ d[918] ^ d[917] ^ d[915] ^ d[909] ^ d[907] ^ d[906] ^ d[905] ^ d[904] ^ d[903] ^ d[900] ^ d[898] ^ d[897] ^ d[894] ^ d[893] ^ d[890] ^ d[888] ^ d[887] ^ d[886] ^ d[884] ^ d[883] ^ d[882] ^ d[881] ^ d[879] ^ d[878] ^ d[875] ^ d[874] ^ d[873] ^ d[870] ^ d[861] ^ d[859] ^ d[857] ^ d[856] ^ d[852] ^ d[851] ^ d[849] ^ d[846] ^ d[843] ^ d[839] ^ d[838] ^ d[837] ^ d[836] ^ d[835] ^ d[832] ^ d[827] ^ d[826] ^ d[825] ^ d[824] ^ d[820] ^ d[816] ^ d[814] ^ d[813] ^ d[812] ^ d[810] ^ d[808] ^ d[807] ^ d[805] ^ d[803] ^ d[801] ^ d[800] ^ d[798] ^ d[797] ^ d[796] ^ d[794] ^ d[791] ^ d[789] ^ d[788] ^ d[787] ^ d[784] ^ d[783] ^ d[782] ^ d[781] ^ d[780] ^ d[775] ^ d[773] ^ d[769] ^ d[768] ^ d[767] ^ d[766] ^ d[765] ^ d[762] ^ d[760] ^ d[759] ^ d[757] ^ d[756] ^ d[749] ^ d[748] ^ d[747] ^ d[746] ^ d[745] ^ d[744] ^ d[742] ^ d[739] ^ d[736] ^ d[735] ^ d[730] ^ d[729] ^ d[728] ^ d[727] ^ d[726] ^ d[725] ^ d[723] ^ d[722] ^ d[721] ^ d[719] ^ d[715] ^ d[714] ^ d[712] ^ d[710] ^ d[709] ^ d[707] ^ d[706] ^ d[704] ^ d[701] ^ d[700] ^ d[697] ^ d[693] ^ d[691] ^ d[690] ^ d[689] ^ d[688] ^ d[686] ^ d[685] ^ d[683] ^ d[681] ^ d[680] ^ d[679] ^ d[674] ^ d[672] ^ d[671] ^ d[670] ^ d[669] ^ d[668] ^ d[667] ^ d[666] ^ d[661] ^ d[660] ^ d[659] ^ d[657] ^ d[656] ^ d[655] ^ d[654] ^ d[653] ^ d[647] ^ d[640] ^ d[639] ^ d[638] ^ d[637] ^ d[634] ^ d[633] ^ d[632] ^ d[631] ^ d[629] ^ d[625] ^ d[623] ^ d[619] ^ d[616] ^ d[615] ^ d[614] ^ d[610] ^ d[605] ^ d[604] ^ d[602] ^ d[597] ^ d[594] ^ d[593] ^ d[590] ^ d[586] ^ d[582] ^ d[581] ^ d[576] ^ d[571] ^ d[569] ^ d[565] ^ d[559] ^ d[557] ^ d[555] ^ d[554] ^ d[552] ^ d[550] ^ d[542] ^ d[541] ^ d[540] ^ d[539] ^ d[537] ^ d[535] ^ d[532] ^ d[529] ^ d[528] ^ d[526] ^ d[523] ^ d[520] ^ d[519] ^ d[518] ^ d[517] ^ d[515] ^ d[511] ^ d[508] ^ d[505] ^ d[504] ^ d[503] ^ d[502] ^ d[501] ^ d[500] ^ d[499] ^ d[498] ^ d[497] ^ d[494] ^ d[492] ^ d[491] ^ d[490] ^ d[489] ^ d[487] ^ d[486] ^ d[485] ^ d[483] ^ d[482] ^ d[479] ^ d[478] ^ d[476] ^ d[474] ^ d[473] ^ d[471] ^ d[468] ^ d[466] ^ d[464] ^ d[460] ^ d[458] ^ d[457] ^ d[456] ^ d[454] ^ d[453] ^ d[452] ^ d[451] ^ d[450] ^ d[449] ^ d[448] ^ d[447] ^ d[444] ^ d[443] ^ d[442] ^ d[438] ^ d[437] ^ d[434] ^ d[432] ^ d[430] ^ d[429] ^ d[428] ^ d[424] ^ d[423] ^ d[421] ^ d[420] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[415] ^ d[412] ^ d[410] ^ d[409] ^ d[407] ^ d[406] ^ d[405] ^ d[404] ^ d[400] ^ d[398] ^ d[397] ^ d[396] ^ d[393] ^ d[390] ^ d[389] ^ d[388] ^ d[386] ^ d[384] ^ d[383] ^ d[382] ^ d[381] ^ d[380] ^ d[379] ^ d[377] ^ d[375] ^ d[374] ^ d[373] ^ d[372] ^ d[371] ^ d[370] ^ d[368] ^ d[367] ^ d[365] ^ d[364] ^ d[363] ^ d[359] ^ d[358] ^ d[357] ^ d[352] ^ d[349] ^ d[348] ^ d[347] ^ d[346] ^ d[345] ^ d[344] ^ d[339] ^ d[337] ^ d[335] ^ d[332] ^ d[331] ^ d[329] ^ d[328] ^ d[326] ^ d[325] ^ d[324] ^ d[323] ^ d[319] ^ d[318] ^ d[317] ^ d[315] ^ d[313] ^ d[312] ^ d[311] ^ d[309] ^ d[307] ^ d[305] ^ d[304] ^ d[299] ^ d[296] ^ d[294] ^ d[292] ^ d[288] ^ d[284] ^ d[282] ^ d[279] ^ d[278] ^ d[277] ^ d[274] ^ d[273] ^ d[272] ^ d[270] ^ d[269] ^ d[264] ^ d[263] ^ d[260] ^ d[259] ^ d[258] ^ d[256] ^ d[255] ^ d[252] ^ d[250] ^ d[247] ^ d[246] ^ d[245] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[234] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[222] ^ d[219] ^ d[216] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[205] ^ d[204] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[195] ^ d[194] ^ d[192] ^ d[186] ^ d[185] ^ d[184] ^ d[178] ^ d[176] ^ d[174] ^ d[172] ^ d[171] ^ d[170] ^ d[168] ^ d[167] ^ d[165] ^ d[164] ^ d[163] ^ d[162] ^ d[160] ^ d[158] ^ d[157] ^ d[155] ^ d[154] ^ d[152] ^ d[145] ^ d[144] ^ d[143] ^ d[141] ^ d[133] ^ d[132] ^ d[131] ^ d[126] ^ d[125] ^ d[119] ^ d[117] ^ d[116] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[103] ^ d[101] ^ d[100] ^ d[98] ^ d[96] ^ d[94] ^ d[93] ^ d[92] ^ d[90] ^ d[89] ^ d[86] ^ d[84] ^ d[79] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[66] ^ d[65] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[54] ^ d[53] ^ d[52] ^ d[47] ^ d[45] ^ d[43] ^ d[42] ^ d[40] ^ d[36] ^ d[33] ^ d[31] ^ d[30] ^ d[29] ^ d[27] ^ d[25] ^ d[24] ^ d[22] ^ d[21] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[10] ^ d[9] ^ d[5] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[9] ^ c[11];
    newcrc[11] = d[1020] ^ d[1018] ^ d[1013] ^ d[1012] ^ d[1010] ^ d[1009] ^ d[1007] ^ d[1006] ^ d[1005] ^ d[998] ^ d[996] ^ d[995] ^ d[993] ^ d[989] ^ d[988] ^ d[986] ^ d[982] ^ d[980] ^ d[979] ^ d[977] ^ d[976] ^ d[975] ^ d[973] ^ d[971] ^ d[970] ^ d[967] ^ d[962] ^ d[960] ^ d[958] ^ d[955] ^ d[954] ^ d[953] ^ d[951] ^ d[949] ^ d[946] ^ d[943] ^ d[935] ^ d[934] ^ d[933] ^ d[931] ^ d[929] ^ d[928] ^ d[927] ^ d[926] ^ d[924] ^ d[919] ^ d[918] ^ d[916] ^ d[910] ^ d[908] ^ d[907] ^ d[906] ^ d[905] ^ d[904] ^ d[901] ^ d[899] ^ d[898] ^ d[895] ^ d[894] ^ d[891] ^ d[889] ^ d[888] ^ d[887] ^ d[885] ^ d[884] ^ d[883] ^ d[882] ^ d[880] ^ d[879] ^ d[876] ^ d[875] ^ d[874] ^ d[871] ^ d[862] ^ d[860] ^ d[858] ^ d[857] ^ d[853] ^ d[852] ^ d[850] ^ d[847] ^ d[844] ^ d[840] ^ d[839] ^ d[838] ^ d[837] ^ d[836] ^ d[833] ^ d[828] ^ d[827] ^ d[826] ^ d[825] ^ d[821] ^ d[817] ^ d[815] ^ d[814] ^ d[813] ^ d[811] ^ d[809] ^ d[808] ^ d[806] ^ d[804] ^ d[802] ^ d[801] ^ d[799] ^ d[798] ^ d[797] ^ d[795] ^ d[792] ^ d[790] ^ d[789] ^ d[788] ^ d[785] ^ d[784] ^ d[783] ^ d[782] ^ d[781] ^ d[776] ^ d[774] ^ d[770] ^ d[769] ^ d[768] ^ d[767] ^ d[766] ^ d[763] ^ d[761] ^ d[760] ^ d[758] ^ d[757] ^ d[750] ^ d[749] ^ d[748] ^ d[747] ^ d[746] ^ d[745] ^ d[743] ^ d[740] ^ d[737] ^ d[736] ^ d[731] ^ d[730] ^ d[729] ^ d[728] ^ d[727] ^ d[726] ^ d[724] ^ d[723] ^ d[722] ^ d[720] ^ d[716] ^ d[715] ^ d[713] ^ d[711] ^ d[710] ^ d[708] ^ d[707] ^ d[705] ^ d[702] ^ d[701] ^ d[698] ^ d[694] ^ d[692] ^ d[691] ^ d[690] ^ d[689] ^ d[687] ^ d[686] ^ d[684] ^ d[682] ^ d[681] ^ d[680] ^ d[675] ^ d[673] ^ d[672] ^ d[671] ^ d[670] ^ d[669] ^ d[668] ^ d[667] ^ d[662] ^ d[661] ^ d[660] ^ d[658] ^ d[657] ^ d[656] ^ d[655] ^ d[654] ^ d[648] ^ d[641] ^ d[640] ^ d[639] ^ d[638] ^ d[635] ^ d[634] ^ d[633] ^ d[632] ^ d[630] ^ d[626] ^ d[624] ^ d[620] ^ d[617] ^ d[616] ^ d[615] ^ d[611] ^ d[606] ^ d[605] ^ d[603] ^ d[598] ^ d[595] ^ d[594] ^ d[591] ^ d[587] ^ d[583] ^ d[582] ^ d[577] ^ d[572] ^ d[570] ^ d[566] ^ d[560] ^ d[558] ^ d[556] ^ d[555] ^ d[553] ^ d[551] ^ d[543] ^ d[542] ^ d[541] ^ d[540] ^ d[538] ^ d[536] ^ d[533] ^ d[530] ^ d[529] ^ d[527] ^ d[524] ^ d[521] ^ d[520] ^ d[519] ^ d[518] ^ d[516] ^ d[512] ^ d[509] ^ d[506] ^ d[505] ^ d[504] ^ d[503] ^ d[502] ^ d[501] ^ d[500] ^ d[499] ^ d[498] ^ d[495] ^ d[493] ^ d[492] ^ d[491] ^ d[490] ^ d[488] ^ d[487] ^ d[486] ^ d[484] ^ d[483] ^ d[480] ^ d[479] ^ d[477] ^ d[475] ^ d[474] ^ d[472] ^ d[469] ^ d[467] ^ d[465] ^ d[461] ^ d[459] ^ d[458] ^ d[457] ^ d[455] ^ d[454] ^ d[453] ^ d[452] ^ d[451] ^ d[450] ^ d[449] ^ d[448] ^ d[445] ^ d[444] ^ d[443] ^ d[439] ^ d[438] ^ d[435] ^ d[433] ^ d[431] ^ d[430] ^ d[429] ^ d[425] ^ d[424] ^ d[422] ^ d[421] ^ d[420] ^ d[419] ^ d[418] ^ d[417] ^ d[416] ^ d[413] ^ d[411] ^ d[410] ^ d[408] ^ d[407] ^ d[406] ^ d[405] ^ d[401] ^ d[399] ^ d[398] ^ d[397] ^ d[394] ^ d[391] ^ d[390] ^ d[389] ^ d[387] ^ d[385] ^ d[384] ^ d[383] ^ d[382] ^ d[381] ^ d[380] ^ d[378] ^ d[376] ^ d[375] ^ d[374] ^ d[373] ^ d[372] ^ d[371] ^ d[369] ^ d[368] ^ d[366] ^ d[365] ^ d[364] ^ d[360] ^ d[359] ^ d[358] ^ d[353] ^ d[350] ^ d[349] ^ d[348] ^ d[347] ^ d[346] ^ d[345] ^ d[340] ^ d[338] ^ d[336] ^ d[333] ^ d[332] ^ d[330] ^ d[329] ^ d[327] ^ d[326] ^ d[325] ^ d[324] ^ d[320] ^ d[319] ^ d[318] ^ d[316] ^ d[314] ^ d[313] ^ d[312] ^ d[310] ^ d[308] ^ d[306] ^ d[305] ^ d[300] ^ d[297] ^ d[295] ^ d[293] ^ d[289] ^ d[285] ^ d[283] ^ d[280] ^ d[279] ^ d[278] ^ d[275] ^ d[274] ^ d[273] ^ d[271] ^ d[270] ^ d[265] ^ d[264] ^ d[261] ^ d[260] ^ d[259] ^ d[257] ^ d[256] ^ d[253] ^ d[251] ^ d[248] ^ d[247] ^ d[246] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[235] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[223] ^ d[220] ^ d[217] ^ d[214] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[206] ^ d[205] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[196] ^ d[195] ^ d[193] ^ d[187] ^ d[186] ^ d[185] ^ d[179] ^ d[177] ^ d[175] ^ d[173] ^ d[172] ^ d[171] ^ d[169] ^ d[168] ^ d[166] ^ d[165] ^ d[164] ^ d[163] ^ d[161] ^ d[159] ^ d[158] ^ d[156] ^ d[155] ^ d[153] ^ d[146] ^ d[145] ^ d[144] ^ d[142] ^ d[134] ^ d[133] ^ d[132] ^ d[127] ^ d[126] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[104] ^ d[102] ^ d[101] ^ d[99] ^ d[97] ^ d[95] ^ d[94] ^ d[93] ^ d[91] ^ d[90] ^ d[87] ^ d[85] ^ d[80] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[67] ^ d[66] ^ d[64] ^ d[63] ^ d[61] ^ d[60] ^ d[59] ^ d[58] ^ d[57] ^ d[55] ^ d[54] ^ d[53] ^ d[48] ^ d[46] ^ d[44] ^ d[43] ^ d[41] ^ d[37] ^ d[34] ^ d[32] ^ d[31] ^ d[30] ^ d[28] ^ d[26] ^ d[25] ^ d[23] ^ d[22] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[14] ^ d[11] ^ d[10] ^ d[6] ^ c[1] ^ c[2] ^ c[4] ^ c[5] ^ c[10] ^ c[12];
    newcrc[12] = d[1023] ^ d[1020] ^ d[1019] ^ d[1017] ^ d[1016] ^ d[1013] ^ d[1012] ^ d[1010] ^ d[1008] ^ d[1007] ^ d[1002] ^ d[998] ^ d[995] ^ d[994] ^ d[993] ^ d[992] ^ d[991] ^ d[989] ^ d[988] ^ d[987] ^ d[986] ^ d[984] ^ d[982] ^ d[980] ^ d[979] ^ d[978] ^ d[977] ^ d[975] ^ d[972] ^ d[971] ^ d[970] ^ d[966] ^ d[964] ^ d[962] ^ d[960] ^ d[959] ^ d[958] ^ d[957] ^ d[956] ^ d[954] ^ d[953] ^ d[951] ^ d[949] ^ d[948] ^ d[947] ^ d[946] ^ d[945] ^ d[944] ^ d[942] ^ d[941] ^ d[938] ^ d[937] ^ d[934] ^ d[933] ^ d[932] ^ d[931] ^ d[929] ^ d[927] ^ d[926] ^ d[924] ^ d[922] ^ d[921] ^ d[920] ^ d[918] ^ d[917] ^ d[915] ^ d[914] ^ d[911] ^ d[910] ^ d[906] ^ d[905] ^ d[904] ^ d[903] ^ d[900] ^ d[899] ^ d[898] ^ d[894] ^ d[892] ^ d[891] ^ d[890] ^ d[887] ^ d[885] ^ d[884] ^ d[883] ^ d[882] ^ d[878] ^ d[877] ^ d[876] ^ d[874] ^ d[871] ^ d[870] ^ d[868] ^ d[867] ^ d[866] ^ d[864] ^ d[863] ^ d[862] ^ d[860] ^ d[858] ^ d[857] ^ d[856] ^ d[855] ^ d[853] ^ d[852] ^ d[851] ^ d[850] ^ d[848] ^ d[846] ^ d[842] ^ d[841] ^ d[838] ^ d[836] ^ d[835] ^ d[833] ^ d[832] ^ d[831] ^ d[830] ^ d[829] ^ d[828] ^ d[827] ^ d[826] ^ d[818] ^ d[812] ^ d[811] ^ d[810] ^ d[807] ^ d[805] ^ d[799] ^ d[798] ^ d[796] ^ d[789] ^ d[787] ^ d[786] ^ d[783] ^ d[781] ^ d[780] ^ d[778] ^ d[777] ^ d[776] ^ d[774] ^ d[772] ^ d[771] ^ d[770] ^ d[768] ^ d[765] ^ d[763] ^ d[761] ^ d[760] ^ d[759] ^ d[758] ^ d[756] ^ d[752] ^ d[748] ^ d[747] ^ d[746] ^ d[745] ^ d[741] ^ d[740] ^ d[736] ^ d[734] ^ d[733] ^ d[732] ^ d[730] ^ d[729] ^ d[727] ^ d[724] ^ d[721] ^ d[719] ^ d[715] ^ d[713] ^ d[712] ^ d[711] ^ d[710] ^ d[709] ^ d[706] ^ d[704] ^ d[700] ^ d[699] ^ d[698] ^ d[696] ^ d[694] ^ d[692] ^ d[691] ^ d[690] ^ d[689] ^ d[685] ^ d[684] ^ d[683] ^ d[680] ^ d[678] ^ d[677] ^ d[676] ^ d[674] ^ d[673] ^ d[668] ^ d[667] ^ d[666] ^ d[665] ^ d[663] ^ d[662] ^ d[661] ^ d[655] ^ d[654] ^ d[653] ^ d[652] ^ d[650] ^ d[649] ^ d[648] ^ d[646] ^ d[644] ^ d[642] ^ d[640] ^ d[637] ^ d[635] ^ d[633] ^ d[632] ^ d[630] ^ d[628] ^ d[627] ^ d[626] ^ d[624] ^ d[622] ^ d[621] ^ d[620] ^ d[618] ^ d[616] ^ d[613] ^ d[609] ^ d[608] ^ d[605] ^ d[604] ^ d[603] ^ d[602] ^ d[601] ^ d[599] ^ d[598] ^ d[597] ^ d[594] ^ d[593] ^ d[592] ^ d[591] ^ d[590] ^ d[589] ^ d[587] ^ d[586] ^ d[585] ^ d[584] ^ d[583] ^ d[582] ^ d[581] ^ d[578] ^ d[577] ^ d[573] ^ d[567] ^ d[557] ^ d[555] ^ d[552] ^ d[551] ^ d[550] ^ d[547] ^ d[546] ^ d[543] ^ d[542] ^ d[540] ^ d[537] ^ d[536] ^ d[535] ^ d[532] ^ d[531] ^ d[530] ^ d[528] ^ d[521] ^ d[518] ^ d[516] ^ d[515] ^ d[514] ^ d[513] ^ d[512] ^ d[511] ^ d[510] ^ d[508] ^ d[507] ^ d[504] ^ d[502] ^ d[501] ^ d[499] ^ d[496] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[486] ^ d[482] ^ d[481] ^ d[480] ^ d[478] ^ d[472] ^ d[471] ^ d[469] ^ d[468] ^ d[467] ^ d[466] ^ d[465] ^ d[463] ^ d[461] ^ d[459] ^ d[458] ^ d[457] ^ d[456] ^ d[453] ^ d[451] ^ d[450] ^ d[448] ^ d[445] ^ d[444] ^ d[442] ^ d[438] ^ d[436] ^ d[435] ^ d[434] ^ d[431] ^ d[428] ^ d[426] ^ d[424] ^ d[421] ^ d[420] ^ d[419] ^ d[418] ^ d[413] ^ d[410] ^ d[409] ^ d[408] ^ d[407] ^ d[406] ^ d[398] ^ d[396] ^ d[395] ^ d[392] ^ d[387] ^ d[386] ^ d[384] ^ d[383] ^ d[381] ^ d[378] ^ d[375] ^ d[374] ^ d[373] ^ d[372] ^ d[366] ^ d[365] ^ d[363] ^ d[359] ^ d[357] ^ d[356] ^ d[353] ^ d[352] ^ d[350] ^ d[349] ^ d[348] ^ d[347] ^ d[342] ^ d[338] ^ d[337] ^ d[335] ^ d[334] ^ d[331] ^ d[329] ^ d[326] ^ d[325] ^ d[324] ^ d[323] ^ d[320] ^ d[319] ^ d[317] ^ d[311] ^ d[310] ^ d[309] ^ d[306] ^ d[303] ^ d[299] ^ d[297] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[291] ^ d[289] ^ d[288] ^ d[287] ^ d[286] ^ d[285] ^ d[284] ^ d[283] ^ d[281] ^ d[279] ^ d[276] ^ d[271] ^ d[270] ^ d[268] ^ d[266] ^ d[264] ^ d[261] ^ d[260] ^ d[258] ^ d[253] ^ d[250] ^ d[249] ^ d[248] ^ d[246] ^ d[243] ^ d[242] ^ d[237] ^ d[236] ^ d[233] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[221] ^ d[219] ^ d[218] ^ d[215] ^ d[210] ^ d[208] ^ d[203] ^ d[202] ^ d[199] ^ d[197] ^ d[196] ^ d[190] ^ d[186] ^ d[184] ^ d[183] ^ d[180] ^ d[179] ^ d[175] ^ d[174] ^ d[172] ^ d[171] ^ d[169] ^ d[167] ^ d[166] ^ d[161] ^ d[160] ^ d[158] ^ d[157] ^ d[155] ^ d[154] ^ d[152] ^ d[151] ^ d[148] ^ d[147] ^ d[144] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[135] ^ d[134] ^ d[133] ^ d[132] ^ d[128] ^ d[123] ^ d[119] ^ d[117] ^ d[114] ^ d[111] ^ d[109] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[100] ^ d[94] ^ d[92] ^ d[91] ^ d[84] ^ d[82] ^ d[80] ^ d[78] ^ d[77] ^ d[76] ^ d[73] ^ d[71] ^ d[70] ^ d[68] ^ d[66] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[59] ^ d[54] ^ d[52] ^ d[51] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[38] ^ d[31] ^ d[29] ^ d[28] ^ d[24] ^ d[23] ^ d[22] ^ d[18] ^ d[16] ^ d[15] ^ d[8] ^ d[7] ^ d[4] ^ d[0] ^ c[0] ^ c[2] ^ c[4] ^ c[5] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[15];
    newcrc[13] = d[1021] ^ d[1020] ^ d[1018] ^ d[1017] ^ d[1014] ^ d[1013] ^ d[1011] ^ d[1009] ^ d[1008] ^ d[1003] ^ d[999] ^ d[996] ^ d[995] ^ d[994] ^ d[993] ^ d[992] ^ d[990] ^ d[989] ^ d[988] ^ d[987] ^ d[985] ^ d[983] ^ d[981] ^ d[980] ^ d[979] ^ d[978] ^ d[976] ^ d[973] ^ d[972] ^ d[971] ^ d[967] ^ d[965] ^ d[963] ^ d[961] ^ d[960] ^ d[959] ^ d[958] ^ d[957] ^ d[955] ^ d[954] ^ d[952] ^ d[950] ^ d[949] ^ d[948] ^ d[947] ^ d[946] ^ d[945] ^ d[943] ^ d[942] ^ d[939] ^ d[938] ^ d[935] ^ d[934] ^ d[933] ^ d[932] ^ d[930] ^ d[928] ^ d[927] ^ d[925] ^ d[923] ^ d[922] ^ d[921] ^ d[919] ^ d[918] ^ d[916] ^ d[915] ^ d[912] ^ d[911] ^ d[907] ^ d[906] ^ d[905] ^ d[904] ^ d[901] ^ d[900] ^ d[899] ^ d[895] ^ d[893] ^ d[892] ^ d[891] ^ d[888] ^ d[886] ^ d[885] ^ d[884] ^ d[883] ^ d[879] ^ d[878] ^ d[877] ^ d[875] ^ d[872] ^ d[871] ^ d[869] ^ d[868] ^ d[867] ^ d[865] ^ d[864] ^ d[863] ^ d[861] ^ d[859] ^ d[858] ^ d[857] ^ d[856] ^ d[854] ^ d[853] ^ d[852] ^ d[851] ^ d[849] ^ d[847] ^ d[843] ^ d[842] ^ d[839] ^ d[837] ^ d[836] ^ d[834] ^ d[833] ^ d[832] ^ d[831] ^ d[830] ^ d[829] ^ d[828] ^ d[827] ^ d[819] ^ d[813] ^ d[812] ^ d[811] ^ d[808] ^ d[806] ^ d[800] ^ d[799] ^ d[797] ^ d[790] ^ d[788] ^ d[787] ^ d[784] ^ d[782] ^ d[781] ^ d[779] ^ d[778] ^ d[777] ^ d[775] ^ d[773] ^ d[772] ^ d[771] ^ d[769] ^ d[766] ^ d[764] ^ d[762] ^ d[761] ^ d[760] ^ d[759] ^ d[757] ^ d[753] ^ d[749] ^ d[748] ^ d[747] ^ d[746] ^ d[742] ^ d[741] ^ d[737] ^ d[735] ^ d[734] ^ d[733] ^ d[731] ^ d[730] ^ d[728] ^ d[725] ^ d[722] ^ d[720] ^ d[716] ^ d[714] ^ d[713] ^ d[712] ^ d[711] ^ d[710] ^ d[707] ^ d[705] ^ d[701] ^ d[700] ^ d[699] ^ d[697] ^ d[695] ^ d[693] ^ d[692] ^ d[691] ^ d[690] ^ d[686] ^ d[685] ^ d[684] ^ d[681] ^ d[679] ^ d[678] ^ d[677] ^ d[675] ^ d[674] ^ d[669] ^ d[668] ^ d[667] ^ d[666] ^ d[664] ^ d[663] ^ d[662] ^ d[656] ^ d[655] ^ d[654] ^ d[653] ^ d[651] ^ d[650] ^ d[649] ^ d[647] ^ d[645] ^ d[643] ^ d[641] ^ d[638] ^ d[636] ^ d[634] ^ d[633] ^ d[631] ^ d[629] ^ d[628] ^ d[627] ^ d[625] ^ d[623] ^ d[622] ^ d[621] ^ d[619] ^ d[617] ^ d[614] ^ d[610] ^ d[609] ^ d[606] ^ d[605] ^ d[604] ^ d[603] ^ d[602] ^ d[600] ^ d[599] ^ d[598] ^ d[595] ^ d[594] ^ d[593] ^ d[592] ^ d[591] ^ d[590] ^ d[588] ^ d[587] ^ d[586] ^ d[585] ^ d[584] ^ d[583] ^ d[582] ^ d[579] ^ d[578] ^ d[574] ^ d[568] ^ d[558] ^ d[556] ^ d[553] ^ d[552] ^ d[551] ^ d[548] ^ d[547] ^ d[544] ^ d[543] ^ d[541] ^ d[538] ^ d[537] ^ d[536] ^ d[533] ^ d[532] ^ d[531] ^ d[529] ^ d[522] ^ d[519] ^ d[517] ^ d[516] ^ d[515] ^ d[514] ^ d[513] ^ d[512] ^ d[511] ^ d[509] ^ d[508] ^ d[505] ^ d[503] ^ d[502] ^ d[500] ^ d[497] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[487] ^ d[483] ^ d[482] ^ d[481] ^ d[479] ^ d[473] ^ d[472] ^ d[470] ^ d[469] ^ d[468] ^ d[467] ^ d[466] ^ d[464] ^ d[462] ^ d[460] ^ d[459] ^ d[458] ^ d[457] ^ d[454] ^ d[452] ^ d[451] ^ d[449] ^ d[446] ^ d[445] ^ d[443] ^ d[439] ^ d[437] ^ d[436] ^ d[435] ^ d[432] ^ d[429] ^ d[427] ^ d[425] ^ d[422] ^ d[421] ^ d[420] ^ d[419] ^ d[414] ^ d[411] ^ d[410] ^ d[409] ^ d[408] ^ d[407] ^ d[399] ^ d[397] ^ d[396] ^ d[393] ^ d[388] ^ d[387] ^ d[385] ^ d[384] ^ d[382] ^ d[379] ^ d[376] ^ d[375] ^ d[374] ^ d[373] ^ d[367] ^ d[366] ^ d[364] ^ d[360] ^ d[358] ^ d[357] ^ d[354] ^ d[353] ^ d[351] ^ d[350] ^ d[349] ^ d[348] ^ d[343] ^ d[339] ^ d[338] ^ d[336] ^ d[335] ^ d[332] ^ d[330] ^ d[327] ^ d[326] ^ d[325] ^ d[324] ^ d[321] ^ d[320] ^ d[318] ^ d[312] ^ d[311] ^ d[310] ^ d[307] ^ d[304] ^ d[300] ^ d[298] ^ d[296] ^ d[295] ^ d[294] ^ d[293] ^ d[292] ^ d[290] ^ d[289] ^ d[288] ^ d[287] ^ d[286] ^ d[285] ^ d[284] ^ d[282] ^ d[280] ^ d[277] ^ d[272] ^ d[271] ^ d[269] ^ d[267] ^ d[265] ^ d[262] ^ d[261] ^ d[259] ^ d[254] ^ d[251] ^ d[250] ^ d[249] ^ d[247] ^ d[244] ^ d[243] ^ d[238] ^ d[237] ^ d[234] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[219] ^ d[216] ^ d[211] ^ d[209] ^ d[204] ^ d[203] ^ d[200] ^ d[198] ^ d[197] ^ d[191] ^ d[187] ^ d[185] ^ d[184] ^ d[181] ^ d[180] ^ d[176] ^ d[175] ^ d[173] ^ d[172] ^ d[170] ^ d[168] ^ d[167] ^ d[162] ^ d[161] ^ d[159] ^ d[158] ^ d[156] ^ d[155] ^ d[153] ^ d[152] ^ d[149] ^ d[148] ^ d[145] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[135] ^ d[134] ^ d[133] ^ d[129] ^ d[124] ^ d[120] ^ d[118] ^ d[115] ^ d[112] ^ d[110] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[101] ^ d[95] ^ d[93] ^ d[92] ^ d[85] ^ d[83] ^ d[81] ^ d[79] ^ d[78] ^ d[77] ^ d[74] ^ d[72] ^ d[71] ^ d[69] ^ d[67] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[55] ^ d[53] ^ d[52] ^ d[49] ^ d[48] ^ d[46] ^ d[45] ^ d[39] ^ d[32] ^ d[30] ^ d[29] ^ d[25] ^ d[24] ^ d[23] ^ d[19] ^ d[17] ^ d[16] ^ d[9] ^ d[8] ^ d[5] ^ d[1] ^ c[0] ^ c[1] ^ c[3] ^ c[5] ^ c[6] ^ c[9] ^ c[10] ^ c[12] ^ c[13];
    newcrc[14] = d[1022] ^ d[1021] ^ d[1019] ^ d[1018] ^ d[1015] ^ d[1014] ^ d[1012] ^ d[1010] ^ d[1009] ^ d[1004] ^ d[1000] ^ d[997] ^ d[996] ^ d[995] ^ d[994] ^ d[993] ^ d[991] ^ d[990] ^ d[989] ^ d[988] ^ d[986] ^ d[984] ^ d[982] ^ d[981] ^ d[980] ^ d[979] ^ d[977] ^ d[974] ^ d[973] ^ d[972] ^ d[968] ^ d[966] ^ d[964] ^ d[962] ^ d[961] ^ d[960] ^ d[959] ^ d[958] ^ d[956] ^ d[955] ^ d[953] ^ d[951] ^ d[950] ^ d[949] ^ d[948] ^ d[947] ^ d[946] ^ d[944] ^ d[943] ^ d[940] ^ d[939] ^ d[936] ^ d[935] ^ d[934] ^ d[933] ^ d[931] ^ d[929] ^ d[928] ^ d[926] ^ d[924] ^ d[923] ^ d[922] ^ d[920] ^ d[919] ^ d[917] ^ d[916] ^ d[913] ^ d[912] ^ d[908] ^ d[907] ^ d[906] ^ d[905] ^ d[902] ^ d[901] ^ d[900] ^ d[896] ^ d[894] ^ d[893] ^ d[892] ^ d[889] ^ d[887] ^ d[886] ^ d[885] ^ d[884] ^ d[880] ^ d[879] ^ d[878] ^ d[876] ^ d[873] ^ d[872] ^ d[870] ^ d[869] ^ d[868] ^ d[866] ^ d[865] ^ d[864] ^ d[862] ^ d[860] ^ d[859] ^ d[858] ^ d[857] ^ d[855] ^ d[854] ^ d[853] ^ d[852] ^ d[850] ^ d[848] ^ d[844] ^ d[843] ^ d[840] ^ d[838] ^ d[837] ^ d[835] ^ d[834] ^ d[833] ^ d[832] ^ d[831] ^ d[830] ^ d[829] ^ d[828] ^ d[820] ^ d[814] ^ d[813] ^ d[812] ^ d[809] ^ d[807] ^ d[801] ^ d[800] ^ d[798] ^ d[791] ^ d[789] ^ d[788] ^ d[785] ^ d[783] ^ d[782] ^ d[780] ^ d[779] ^ d[778] ^ d[776] ^ d[774] ^ d[773] ^ d[772] ^ d[770] ^ d[767] ^ d[765] ^ d[763] ^ d[762] ^ d[761] ^ d[760] ^ d[758] ^ d[754] ^ d[750] ^ d[749] ^ d[748] ^ d[747] ^ d[743] ^ d[742] ^ d[738] ^ d[736] ^ d[735] ^ d[734] ^ d[732] ^ d[731] ^ d[729] ^ d[726] ^ d[723] ^ d[721] ^ d[717] ^ d[715] ^ d[714] ^ d[713] ^ d[712] ^ d[711] ^ d[708] ^ d[706] ^ d[702] ^ d[701] ^ d[700] ^ d[698] ^ d[696] ^ d[694] ^ d[693] ^ d[692] ^ d[691] ^ d[687] ^ d[686] ^ d[685] ^ d[682] ^ d[680] ^ d[679] ^ d[678] ^ d[676] ^ d[675] ^ d[670] ^ d[669] ^ d[668] ^ d[667] ^ d[665] ^ d[664] ^ d[663] ^ d[657] ^ d[656] ^ d[655] ^ d[654] ^ d[652] ^ d[651] ^ d[650] ^ d[648] ^ d[646] ^ d[644] ^ d[642] ^ d[639] ^ d[637] ^ d[635] ^ d[634] ^ d[632] ^ d[630] ^ d[629] ^ d[628] ^ d[626] ^ d[624] ^ d[623] ^ d[622] ^ d[620] ^ d[618] ^ d[615] ^ d[611] ^ d[610] ^ d[607] ^ d[606] ^ d[605] ^ d[604] ^ d[603] ^ d[601] ^ d[600] ^ d[599] ^ d[596] ^ d[595] ^ d[594] ^ d[593] ^ d[592] ^ d[591] ^ d[589] ^ d[588] ^ d[587] ^ d[586] ^ d[585] ^ d[584] ^ d[583] ^ d[580] ^ d[579] ^ d[575] ^ d[569] ^ d[559] ^ d[557] ^ d[554] ^ d[553] ^ d[552] ^ d[549] ^ d[548] ^ d[545] ^ d[544] ^ d[542] ^ d[539] ^ d[538] ^ d[537] ^ d[534] ^ d[533] ^ d[532] ^ d[530] ^ d[523] ^ d[520] ^ d[518] ^ d[517] ^ d[516] ^ d[515] ^ d[514] ^ d[513] ^ d[512] ^ d[510] ^ d[509] ^ d[506] ^ d[504] ^ d[503] ^ d[501] ^ d[498] ^ d[492] ^ d[491] ^ d[490] ^ d[489] ^ d[488] ^ d[484] ^ d[483] ^ d[482] ^ d[480] ^ d[474] ^ d[473] ^ d[471] ^ d[470] ^ d[469] ^ d[468] ^ d[467] ^ d[465] ^ d[463] ^ d[461] ^ d[460] ^ d[459] ^ d[458] ^ d[455] ^ d[453] ^ d[452] ^ d[450] ^ d[447] ^ d[446] ^ d[444] ^ d[440] ^ d[438] ^ d[437] ^ d[436] ^ d[433] ^ d[430] ^ d[428] ^ d[426] ^ d[423] ^ d[422] ^ d[421] ^ d[420] ^ d[415] ^ d[412] ^ d[411] ^ d[410] ^ d[409] ^ d[408] ^ d[400] ^ d[398] ^ d[397] ^ d[394] ^ d[389] ^ d[388] ^ d[386] ^ d[385] ^ d[383] ^ d[380] ^ d[377] ^ d[376] ^ d[375] ^ d[374] ^ d[368] ^ d[367] ^ d[365] ^ d[361] ^ d[359] ^ d[358] ^ d[355] ^ d[354] ^ d[352] ^ d[351] ^ d[350] ^ d[349] ^ d[344] ^ d[340] ^ d[339] ^ d[337] ^ d[336] ^ d[333] ^ d[331] ^ d[328] ^ d[327] ^ d[326] ^ d[325] ^ d[322] ^ d[321] ^ d[319] ^ d[313] ^ d[312] ^ d[311] ^ d[308] ^ d[305] ^ d[301] ^ d[299] ^ d[297] ^ d[296] ^ d[295] ^ d[294] ^ d[293] ^ d[291] ^ d[290] ^ d[289] ^ d[288] ^ d[287] ^ d[286] ^ d[285] ^ d[283] ^ d[281] ^ d[278] ^ d[273] ^ d[272] ^ d[270] ^ d[268] ^ d[266] ^ d[263] ^ d[262] ^ d[260] ^ d[255] ^ d[252] ^ d[251] ^ d[250] ^ d[248] ^ d[245] ^ d[244] ^ d[239] ^ d[238] ^ d[235] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[221] ^ d[220] ^ d[217] ^ d[212] ^ d[210] ^ d[205] ^ d[204] ^ d[201] ^ d[199] ^ d[198] ^ d[192] ^ d[188] ^ d[186] ^ d[185] ^ d[182] ^ d[181] ^ d[177] ^ d[176] ^ d[174] ^ d[173] ^ d[171] ^ d[169] ^ d[168] ^ d[163] ^ d[162] ^ d[160] ^ d[159] ^ d[157] ^ d[156] ^ d[154] ^ d[153] ^ d[150] ^ d[149] ^ d[146] ^ d[144] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[135] ^ d[134] ^ d[130] ^ d[125] ^ d[121] ^ d[119] ^ d[116] ^ d[113] ^ d[111] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[102] ^ d[96] ^ d[94] ^ d[93] ^ d[86] ^ d[84] ^ d[82] ^ d[80] ^ d[79] ^ d[78] ^ d[75] ^ d[73] ^ d[72] ^ d[70] ^ d[68] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[56] ^ d[54] ^ d[53] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[40] ^ d[33] ^ d[31] ^ d[30] ^ d[26] ^ d[25] ^ d[24] ^ d[20] ^ d[18] ^ d[17] ^ d[10] ^ d[9] ^ d[6] ^ d[2] ^ c[1] ^ c[2] ^ c[4] ^ c[6] ^ c[7] ^ c[10] ^ c[11] ^ c[13] ^ c[14];
    newcrc[15] = d[1023] ^ d[1022] ^ d[1020] ^ d[1019] ^ d[1016] ^ d[1015] ^ d[1013] ^ d[1011] ^ d[1010] ^ d[1005] ^ d[1001] ^ d[998] ^ d[997] ^ d[996] ^ d[995] ^ d[994] ^ d[992] ^ d[991] ^ d[990] ^ d[989] ^ d[987] ^ d[985] ^ d[983] ^ d[982] ^ d[981] ^ d[980] ^ d[978] ^ d[975] ^ d[974] ^ d[973] ^ d[969] ^ d[967] ^ d[965] ^ d[963] ^ d[962] ^ d[961] ^ d[960] ^ d[959] ^ d[957] ^ d[956] ^ d[954] ^ d[952] ^ d[951] ^ d[950] ^ d[949] ^ d[948] ^ d[947] ^ d[945] ^ d[944] ^ d[941] ^ d[940] ^ d[937] ^ d[936] ^ d[935] ^ d[934] ^ d[932] ^ d[930] ^ d[929] ^ d[927] ^ d[925] ^ d[924] ^ d[923] ^ d[921] ^ d[920] ^ d[918] ^ d[917] ^ d[914] ^ d[913] ^ d[909] ^ d[908] ^ d[907] ^ d[906] ^ d[903] ^ d[902] ^ d[901] ^ d[897] ^ d[895] ^ d[894] ^ d[893] ^ d[890] ^ d[888] ^ d[887] ^ d[886] ^ d[885] ^ d[881] ^ d[880] ^ d[879] ^ d[877] ^ d[874] ^ d[873] ^ d[871] ^ d[870] ^ d[869] ^ d[867] ^ d[866] ^ d[865] ^ d[863] ^ d[861] ^ d[860] ^ d[859] ^ d[858] ^ d[856] ^ d[855] ^ d[854] ^ d[853] ^ d[851] ^ d[849] ^ d[845] ^ d[844] ^ d[841] ^ d[839] ^ d[838] ^ d[836] ^ d[835] ^ d[834] ^ d[833] ^ d[832] ^ d[831] ^ d[830] ^ d[829] ^ d[821] ^ d[815] ^ d[814] ^ d[813] ^ d[810] ^ d[808] ^ d[802] ^ d[801] ^ d[799] ^ d[792] ^ d[790] ^ d[789] ^ d[786] ^ d[784] ^ d[783] ^ d[781] ^ d[780] ^ d[779] ^ d[777] ^ d[775] ^ d[774] ^ d[773] ^ d[771] ^ d[768] ^ d[766] ^ d[764] ^ d[763] ^ d[762] ^ d[761] ^ d[759] ^ d[755] ^ d[751] ^ d[750] ^ d[749] ^ d[748] ^ d[744] ^ d[743] ^ d[739] ^ d[737] ^ d[736] ^ d[735] ^ d[733] ^ d[732] ^ d[730] ^ d[727] ^ d[724] ^ d[722] ^ d[718] ^ d[716] ^ d[715] ^ d[714] ^ d[713] ^ d[712] ^ d[709] ^ d[707] ^ d[703] ^ d[702] ^ d[701] ^ d[699] ^ d[697] ^ d[695] ^ d[694] ^ d[693] ^ d[692] ^ d[688] ^ d[687] ^ d[686] ^ d[683] ^ d[681] ^ d[680] ^ d[679] ^ d[677] ^ d[676] ^ d[671] ^ d[670] ^ d[669] ^ d[668] ^ d[666] ^ d[665] ^ d[664] ^ d[658] ^ d[657] ^ d[656] ^ d[655] ^ d[653] ^ d[652] ^ d[651] ^ d[649] ^ d[647] ^ d[645] ^ d[643] ^ d[640] ^ d[638] ^ d[636] ^ d[635] ^ d[633] ^ d[631] ^ d[630] ^ d[629] ^ d[627] ^ d[625] ^ d[624] ^ d[623] ^ d[621] ^ d[619] ^ d[616] ^ d[612] ^ d[611] ^ d[608] ^ d[607] ^ d[606] ^ d[605] ^ d[604] ^ d[602] ^ d[601] ^ d[600] ^ d[597] ^ d[596] ^ d[595] ^ d[594] ^ d[593] ^ d[592] ^ d[590] ^ d[589] ^ d[588] ^ d[587] ^ d[586] ^ d[585] ^ d[584] ^ d[581] ^ d[580] ^ d[576] ^ d[570] ^ d[560] ^ d[558] ^ d[555] ^ d[554] ^ d[553] ^ d[550] ^ d[549] ^ d[546] ^ d[545] ^ d[543] ^ d[540] ^ d[539] ^ d[538] ^ d[535] ^ d[534] ^ d[533] ^ d[531] ^ d[524] ^ d[521] ^ d[519] ^ d[518] ^ d[517] ^ d[516] ^ d[515] ^ d[514] ^ d[513] ^ d[511] ^ d[510] ^ d[507] ^ d[505] ^ d[504] ^ d[502] ^ d[499] ^ d[493] ^ d[492] ^ d[491] ^ d[490] ^ d[489] ^ d[485] ^ d[484] ^ d[483] ^ d[481] ^ d[475] ^ d[474] ^ d[472] ^ d[471] ^ d[470] ^ d[469] ^ d[468] ^ d[466] ^ d[464] ^ d[462] ^ d[461] ^ d[460] ^ d[459] ^ d[456] ^ d[454] ^ d[453] ^ d[451] ^ d[448] ^ d[447] ^ d[445] ^ d[441] ^ d[439] ^ d[438] ^ d[437] ^ d[434] ^ d[431] ^ d[429] ^ d[427] ^ d[424] ^ d[423] ^ d[422] ^ d[421] ^ d[416] ^ d[413] ^ d[412] ^ d[411] ^ d[410] ^ d[409] ^ d[401] ^ d[399] ^ d[398] ^ d[395] ^ d[390] ^ d[389] ^ d[387] ^ d[386] ^ d[384] ^ d[381] ^ d[378] ^ d[377] ^ d[376] ^ d[375] ^ d[369] ^ d[368] ^ d[366] ^ d[362] ^ d[360] ^ d[359] ^ d[356] ^ d[355] ^ d[353] ^ d[352] ^ d[351] ^ d[350] ^ d[345] ^ d[341] ^ d[340] ^ d[338] ^ d[337] ^ d[334] ^ d[332] ^ d[329] ^ d[328] ^ d[327] ^ d[326] ^ d[323] ^ d[322] ^ d[320] ^ d[314] ^ d[313] ^ d[312] ^ d[309] ^ d[306] ^ d[302] ^ d[300] ^ d[298] ^ d[297] ^ d[296] ^ d[295] ^ d[294] ^ d[292] ^ d[291] ^ d[290] ^ d[289] ^ d[288] ^ d[287] ^ d[286] ^ d[284] ^ d[282] ^ d[279] ^ d[274] ^ d[273] ^ d[271] ^ d[269] ^ d[267] ^ d[264] ^ d[263] ^ d[261] ^ d[256] ^ d[253] ^ d[252] ^ d[251] ^ d[249] ^ d[246] ^ d[245] ^ d[240] ^ d[239] ^ d[236] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[222] ^ d[221] ^ d[218] ^ d[213] ^ d[211] ^ d[206] ^ d[205] ^ d[202] ^ d[200] ^ d[199] ^ d[193] ^ d[189] ^ d[187] ^ d[186] ^ d[183] ^ d[182] ^ d[178] ^ d[177] ^ d[175] ^ d[174] ^ d[172] ^ d[170] ^ d[169] ^ d[164] ^ d[163] ^ d[161] ^ d[160] ^ d[158] ^ d[157] ^ d[155] ^ d[154] ^ d[151] ^ d[150] ^ d[147] ^ d[145] ^ d[144] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[135] ^ d[131] ^ d[126] ^ d[122] ^ d[120] ^ d[117] ^ d[114] ^ d[112] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[103] ^ d[97] ^ d[95] ^ d[94] ^ d[87] ^ d[85] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[76] ^ d[74] ^ d[73] ^ d[71] ^ d[69] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[57] ^ d[55] ^ d[54] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[41] ^ d[34] ^ d[32] ^ d[31] ^ d[27] ^ d[26] ^ d[25] ^ d[21] ^ d[19] ^ d[18] ^ d[11] ^ d[10] ^ d[7] ^ d[3] ^ c[2] ^ c[3] ^ c[5] ^ c[7] ^ c[8] ^ c[11] ^ c[12] ^ c[14] ^ c[15];
    nextCRC16_D1024 = newcrc;
  end
  
endmodule
