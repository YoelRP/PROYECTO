module inv(
  in
  out   );
    output reg  out;
    input wire in ;
assign out = ~in ;

endmodule